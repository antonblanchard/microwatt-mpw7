* NGSPICE file created from multiply_add_64x64.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fa_2 abstract view
.subckt sky130_fd_sc_hd__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fa_1 abstract view
.subckt sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ha_1 abstract view
.subckt sky130_fd_sc_hd__ha_1 A B VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ha_2 abstract view
.subckt sky130_fd_sc_hd__ha_2 A B VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ha_4 abstract view
.subckt sky130_fd_sc_hd__ha_4 A B VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

.subckt multiply_add_64x64 VGND VPWR a[0] a[10] a[11] a[12] a[13] a[14] a[15] a[16]
+ a[17] a[18] a[19] a[1] a[20] a[21] a[22] a[23] a[24] a[25] a[26] a[27] a[28] a[29]
+ a[2] a[30] a[31] a[32] a[33] a[34] a[35] a[36] a[37] a[38] a[39] a[3] a[40] a[41]
+ a[42] a[43] a[44] a[45] a[46] a[47] a[48] a[49] a[4] a[50] a[51] a[52] a[53] a[54]
+ a[55] a[56] a[57] a[58] a[59] a[5] a[60] a[61] a[62] a[63] a[6] a[7] a[8] a[9] b[0]
+ b[10] b[11] b[12] b[13] b[14] b[15] b[16] b[17] b[18] b[19] b[1] b[20] b[21] b[22]
+ b[23] b[24] b[25] b[26] b[27] b[28] b[29] b[2] b[30] b[31] b[32] b[33] b[34] b[35]
+ b[36] b[37] b[38] b[39] b[3] b[40] b[41] b[42] b[43] b[44] b[45] b[46] b[47] b[48]
+ b[49] b[4] b[50] b[51] b[52] b[53] b[54] b[55] b[56] b[57] b[58] b[59] b[5] b[60]
+ b[61] b[62] b[63] b[6] b[7] b[8] b[9] c[0] c[100] c[101] c[102] c[103] c[104] c[105]
+ c[106] c[107] c[108] c[109] c[10] c[110] c[111] c[112] c[113] c[114] c[115] c[116]
+ c[117] c[118] c[119] c[11] c[120] c[121] c[122] c[123] c[124] c[125] c[126] c[127]
+ c[12] c[13] c[14] c[15] c[16] c[17] c[18] c[19] c[1] c[20] c[21] c[22] c[23] c[24]
+ c[25] c[26] c[27] c[28] c[29] c[2] c[30] c[31] c[32] c[33] c[34] c[35] c[36] c[37]
+ c[38] c[39] c[3] c[40] c[41] c[42] c[43] c[44] c[45] c[46] c[47] c[48] c[49] c[4]
+ c[50] c[51] c[52] c[53] c[54] c[55] c[56] c[57] c[58] c[59] c[5] c[60] c[61] c[62]
+ c[63] c[64] c[65] c[66] c[67] c[68] c[69] c[6] c[70] c[71] c[72] c[73] c[74] c[75]
+ c[76] c[77] c[78] c[79] c[7] c[80] c[81] c[82] c[83] c[84] c[85] c[86] c[87] c[88]
+ c[89] c[8] c[90] c[91] c[92] c[93] c[94] c[95] c[96] c[97] c[98] c[99] c[9] clk
+ o[0] o[100] o[101] o[102] o[103] o[104] o[105] o[106] o[107] o[108] o[109] o[10]
+ o[110] o[111] o[112] o[113] o[114] o[115] o[116] o[117] o[118] o[119] o[11] o[120]
+ o[121] o[122] o[123] o[124] o[125] o[126] o[127] o[12] o[13] o[14] o[15] o[16] o[17]
+ o[18] o[19] o[1] o[20] o[21] o[22] o[23] o[24] o[25] o[26] o[27] o[28] o[29] o[2]
+ o[30] o[31] o[32] o[33] o[34] o[35] o[36] o[37] o[38] o[39] o[3] o[40] o[41] o[42]
+ o[43] o[44] o[45] o[46] o[47] o[48] o[49] o[4] o[50] o[51] o[52] o[53] o[54] o[55]
+ o[56] o[57] o[58] o[59] o[5] o[60] o[61] o[62] o[63] o[64] o[65] o[66] o[67] o[68]
+ o[69] o[6] o[70] o[71] o[72] o[73] o[74] o[75] o[76] o[77] o[78] o[79] o[7] o[80]
+ o[81] o[82] o[83] o[84] o[85] o[86] o[87] o[88] o[89] o[8] o[90] o[91] o[92] o[93]
+ o[94] o[95] o[96] o[97] o[98] o[99] o[9] rst
XFILLER_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_57_8 dadda_fa_1_57_8/A dadda_fa_1_57_8/B dadda_fa_1_57_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_58_3/A dadda_fa_3_57_0/A sky130_fd_sc_hd__fa_2
XFILLER_94_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_104_0 dadda_fa_2_104_0/A U$$2875/X U$$3008/X VGND VGND VPWR VPWR dadda_fa_3_105_2/CIN
+ dadda_fa_3_104_3/B sky130_fd_sc_hd__fa_1
XFILLER_74_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1290 U$$1290/A U$$1294/B VGND VGND VPWR VPWR U$$1290/X sky130_fd_sc_hd__xor2_1
XFILLER_167_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_90_2 U$$2581/X U$$2714/X U$$2847/X VGND VGND VPWR VPWR dadda_fa_2_91_4/CIN
+ dadda_fa_2_90_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4513_1904 VGND VGND VPWR VPWR U$$4513_1904/HI U$$4513/B sky130_fd_sc_hd__conb_1
Xdadda_fa_1_83_1 U$$1769/X U$$1902/X U$$2035/X VGND VGND VPWR VPWR dadda_fa_2_84_2/A
+ dadda_fa_2_83_4/B sky130_fd_sc_hd__fa_1
XFILLER_104_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_60_0 dadda_fa_4_60_0/A dadda_fa_4_60_0/B dadda_fa_4_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_61_0/A dadda_fa_5_60_1/A sky130_fd_sc_hd__fa_1
Xfanout820 U$$2471/X VGND VGND VPWR VPWR fanout820/X sky130_fd_sc_hd__clkbuf_16
XFILLER_132_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_76_0 U$$1489/X U$$1622/X U$$1755/X VGND VGND VPWR VPWR dadda_fa_2_77_0/B
+ dadda_fa_2_76_3/B sky130_fd_sc_hd__fa_1
Xfanout831 U$$2282/B2 VGND VGND VPWR VPWR U$$2252/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_120_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout842 U$$2181/B2 VGND VGND VPWR VPWR U$$2189/B2 sky130_fd_sc_hd__buf_6
Xfanout853 U$$1859/B2 VGND VGND VPWR VPWR U$$1829/B2 sky130_fd_sc_hd__buf_4
XFILLER_131_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout864 U$$1760/B2 VGND VGND VPWR VPWR U$$1726/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout875 U$$1621/B2 VGND VGND VPWR VPWR U$$1587/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout886 U$$253/B2 VGND VGND VPWR VPWR U$$207/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout897 U$$1361/B2 VGND VGND VPWR VPWR U$$1327/B2 sky130_fd_sc_hd__buf_4
XFILLER_58_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3609 U$$3609/A U$$3615/B VGND VGND VPWR VPWR U$$3609/X sky130_fd_sc_hd__xor2_1
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2908 U$$2908/A U$$2944/B VGND VGND VPWR VPWR U$$2908/X sky130_fd_sc_hd__xor2_1
XU$$2919 U$$999/B1 U$$2937/A2 U$$866/A1 U$$2937/B2 VGND VGND VPWR VPWR U$$2920/A sky130_fd_sc_hd__a22o_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_5_124_1 U$$4511/X input156/X VGND VGND VPWR VPWR dadda_fa_6_125_0/CIN dadda_fa_7_124_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_363_ _364_/CLK _363_/D VGND VGND VPWR VPWR _363_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_294_ _422_/CLK _294_/D VGND VGND VPWR VPWR _294_/Q sky130_fd_sc_hd__dfxtp_1
XU$$3431_1820 VGND VGND VPWR VPWR U$$3431_1820/HI U$$3431/A1 sky130_fd_sc_hd__conb_1
XFILLER_6_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_98_1 dadda_fa_3_98_1/A dadda_fa_3_98_1/B dadda_fa_3_98_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_99_0/CIN dadda_fa_4_98_2/A sky130_fd_sc_hd__fa_1
XFILLER_6_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_75_0 dadda_fa_6_75_0/A dadda_fa_6_75_0/B dadda_fa_6_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_76_0/B dadda_fa_7_75_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_174_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_915 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$370 U$$505/B1 U$$408/A2 U$$370/B1 U$$408/B2 VGND VGND VPWR VPWR U$$371/A sky130_fd_sc_hd__a22o_1
XFILLER_91_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$381 U$$381/A U$$387/B VGND VGND VPWR VPWR U$$381/X sky130_fd_sc_hd__xor2_1
XU$$392 U$$940/A1 U$$408/A2 U$$942/A1 U$$408/B2 VGND VGND VPWR VPWR U$$393/A sky130_fd_sc_hd__a22o_1
XFILLER_33_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_93_0 U$$2853/X U$$2986/X U$$3119/X VGND VGND VPWR VPWR dadda_fa_3_94_0/B
+ dadda_fa_3_93_2/B sky130_fd_sc_hd__fa_1
XFILLER_173_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_62_6 dadda_fa_1_62_6/A dadda_fa_1_62_6/B dadda_fa_1_62_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_63_2/B dadda_fa_2_62_5/B sky130_fd_sc_hd__fa_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_55_5 U$$2777/X U$$2910/X U$$3043/X VGND VGND VPWR VPWR dadda_fa_2_56_2/A
+ dadda_fa_2_55_5/A sky130_fd_sc_hd__fa_1
XFILLER_95_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_48_4 U$$1699/X U$$1832/X U$$1965/X VGND VGND VPWR VPWR dadda_fa_2_49_2/B
+ dadda_fa_2_48_5/A sky130_fd_sc_hd__fa_1
XFILLER_103_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_18_2 dadda_fa_4_18_2/A dadda_fa_4_18_2/B dadda_ha_3_18_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_19_0/CIN dadda_fa_5_18_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_92_0 dadda_fa_7_92_0/A dadda_fa_7_92_0/B dadda_fa_7_92_0/CIN VGND VGND
+ VPWR VPWR _389_/D _260_/D sky130_fd_sc_hd__fa_2
XFILLER_164_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1604 U$$2862/B1 VGND VGND VPWR VPWR U$$946/A1 sky130_fd_sc_hd__buf_4
Xfanout1615 U$$4506/A1 VGND VGND VPWR VPWR U$$3684/A1 sky130_fd_sc_hd__buf_4
XFILLER_132_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1626 U$$2860/A1 VGND VGND VPWR VPWR U$$4504/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1637 U$$938/A1 VGND VGND VPWR VPWR U$$936/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_104_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout650 U$$1218/A2 VGND VGND VPWR VPWR U$$1226/A2 sky130_fd_sc_hd__buf_6
Xfanout1648 U$$2578/B1 VGND VGND VPWR VPWR U$$386/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout661 U$$952/B2 VGND VGND VPWR VPWR U$$902/B2 sky130_fd_sc_hd__clkbuf_8
XU$$4107 U$$4107/A1 U$$4107/A2 U$$4107/B1 U$$4107/B2 VGND VGND VPWR VPWR U$$4108/A
+ sky130_fd_sc_hd__a22o_1
XU$$3422_1819 VGND VGND VPWR VPWR U$$3422_1819/HI U$$3422/B1 sky130_fd_sc_hd__conb_1
Xfanout1659 U$$4496/A1 VGND VGND VPWR VPWR U$$4220/B1 sky130_fd_sc_hd__buf_4
XU$$4118 U$$4392/A1 U$$4158/A2 U$$4257/A1 U$$4158/B2 VGND VGND VPWR VPWR U$$4119/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout672 U$$771/B2 VGND VGND VPWR VPWR U$$743/B2 sky130_fd_sc_hd__clkbuf_4
XU$$4129 U$$4129/A U$$4133/B VGND VGND VPWR VPWR U$$4129/X sky130_fd_sc_hd__xor2_1
XFILLER_77_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout683 U$$553/X VGND VGND VPWR VPWR U$$642/B2 sky130_fd_sc_hd__buf_4
Xfanout694 U$$543/B2 VGND VGND VPWR VPWR U$$501/B2 sky130_fd_sc_hd__buf_4
XFILLER_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3406 U$$4226/B1 U$$3416/A2 U$$4093/A1 U$$3416/B2 VGND VGND VPWR VPWR U$$3407/A
+ sky130_fd_sc_hd__a22o_1
XU$$3417 U$$3417/A U$$3417/B VGND VGND VPWR VPWR U$$3417/X sky130_fd_sc_hd__xor2_1
XU$$3428 U$$3562/A U$$3428/B VGND VGND VPWR VPWR U$$3428/X sky130_fd_sc_hd__and2_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3439 U$$3713/A1 U$$3439/A2 U$$3713/B1 U$$3439/B2 VGND VGND VPWR VPWR U$$3440/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_160_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2705 U$$2840/B1 U$$2707/A2 U$$2707/A1 U$$2707/B2 VGND VGND VPWR VPWR U$$2706/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2716 U$$2716/A U$$2739/A VGND VGND VPWR VPWR U$$2716/X sky130_fd_sc_hd__xor2_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2727 U$$946/A1 U$$2737/A2 U$$948/A1 U$$2737/B2 VGND VGND VPWR VPWR U$$2728/A sky130_fd_sc_hd__a22o_1
XFILLER_37_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2738 U$$2738/A U$$2738/B VGND VGND VPWR VPWR U$$2738/X sky130_fd_sc_hd__xor2_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2749 U$$2749/A U$$2805/B VGND VGND VPWR VPWR U$$2749/X sky130_fd_sc_hd__xor2_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_2 U$$845/X U$$978/X U$$1111/X VGND VGND VPWR VPWR dadda_fa_4_21_1/A
+ dadda_fa_4_20_2/B sky130_fd_sc_hd__fa_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_415_ _415_/CLK _415_/D VGND VGND VPWR VPWR _415_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_346_ _346_/CLK _346_/D VGND VGND VPWR VPWR _346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_277_ _405_/CLK _277_/D VGND VGND VPWR VPWR _277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_72_5 dadda_fa_2_72_5/A dadda_fa_2_72_5/B dadda_fa_2_72_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_2/A dadda_fa_4_72_0/A sky130_fd_sc_hd__fa_1
XFILLER_97_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_65_4 dadda_fa_2_65_4/A dadda_fa_2_65_4/B dadda_fa_2_65_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_1/CIN dadda_fa_3_65_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_110_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_58_3 dadda_fa_2_58_3/A dadda_fa_2_58_3/B dadda_fa_2_58_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_1/B dadda_fa_3_58_3/B sky130_fd_sc_hd__fa_1
Xdadda_fa_5_28_1 dadda_fa_5_28_1/A dadda_fa_5_28_1/B dadda_fa_5_28_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_29_0/B dadda_fa_7_28_0/A sky130_fd_sc_hd__fa_2
XU$$3940 U$$4488/A1 U$$3948/A2 U$$4490/A1 U$$3948/B2 VGND VGND VPWR VPWR U$$3941/A
+ sky130_fd_sc_hd__a22o_1
XU$$3951 U$$3951/A U$$3965/B VGND VGND VPWR VPWR U$$3951/X sky130_fd_sc_hd__xor2_1
XFILLER_25_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3962 U$$4508/B1 U$$3970/A2 U$$3964/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3963/A
+ sky130_fd_sc_hd__a22o_1
XU$$3973 U$$3973/A VGND VGND VPWR VPWR U$$3973/Y sky130_fd_sc_hd__inv_1
XFILLER_18_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3984 U$$3984/A U$$4026/B VGND VGND VPWR VPWR U$$3984/X sky130_fd_sc_hd__xor2_1
XU$$3995 U$$4132/A1 U$$4025/A2 U$$4132/B1 U$$4025/B2 VGND VGND VPWR VPWR U$$3996/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_102_1 dadda_fa_5_102_1/A dadda_fa_5_102_1/B dadda_fa_5_102_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_103_0/B dadda_fa_7_102_0/A sky130_fd_sc_hd__fa_1
XFILLER_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput264 output264/A VGND VGND VPWR VPWR o[106] sky130_fd_sc_hd__buf_2
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput275 output275/A VGND VGND VPWR VPWR o[116] sky130_fd_sc_hd__buf_2
Xoutput286 output286/A VGND VGND VPWR VPWR o[126] sky130_fd_sc_hd__buf_2
XFILLER_87_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput297 output297/A VGND VGND VPWR VPWR o[20] sky130_fd_sc_hd__buf_2
XU$$2061_1798 VGND VGND VPWR VPWR U$$2061_1798/HI U$$2061/A1 sky130_fd_sc_hd__conb_1
XFILLER_87_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_60_3 U$$3186/X U$$3319/X U$$3452/X VGND VGND VPWR VPWR dadda_fa_2_61_1/B
+ dadda_fa_2_60_4/B sky130_fd_sc_hd__fa_1
XFILLER_114_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_2 U$$1177/X U$$1310/X U$$1443/X VGND VGND VPWR VPWR dadda_fa_2_54_1/A
+ dadda_fa_2_53_4/A sky130_fd_sc_hd__fa_1
XFILLER_56_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_30_1 dadda_fa_4_30_1/A dadda_fa_4_30_1/B dadda_fa_4_30_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_31_0/B dadda_fa_5_30_1/B sky130_fd_sc_hd__fa_1
XFILLER_28_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_46_1 U$$498/X U$$631/X U$$764/X VGND VGND VPWR VPWR dadda_fa_2_47_2/A
+ dadda_fa_2_46_4/B sky130_fd_sc_hd__fa_1
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_23_0 dadda_fa_4_23_0/A dadda_fa_4_23_0/B dadda_fa_4_23_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_24_0/A dadda_fa_5_23_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_39_0 U$$85/X U$$218/X U$$351/X VGND VGND VPWR VPWR dadda_fa_2_40_4/A dadda_fa_2_39_5/B
+ sky130_fd_sc_hd__fa_1
XFILLER_82_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_200_ _328_/CLK _200_/D VGND VGND VPWR VPWR _200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1105 final_adder.U$$174/B final_adder.U$$945/X VGND VGND VPWR VPWR
+ output364/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1116 final_adder.U$$162/A final_adder.U$$871/X VGND VGND VPWR VPWR
+ output376/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1127 final_adder.U$$152/B final_adder.U$$923/X VGND VGND VPWR VPWR
+ output261/A sky130_fd_sc_hd__xor2_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1138 final_adder.U$$140/A final_adder.U$$849/X VGND VGND VPWR VPWR
+ output273/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1149 final_adder.U$$130/B final_adder.U$$901/X VGND VGND VPWR VPWR
+ output285/A sky130_fd_sc_hd__xor2_1
XFILLER_137_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_75_3 dadda_fa_3_75_3/A dadda_fa_3_75_3/B dadda_fa_3_75_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_1/B dadda_fa_4_75_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_133_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1401 input34/X VGND VGND VPWR VPWR U$$254/B sky130_fd_sc_hd__buf_6
Xdadda_fa_3_68_2 dadda_fa_3_68_2/A dadda_fa_3_68_2/B dadda_fa_3_68_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_1/A dadda_fa_4_68_2/B sky130_fd_sc_hd__fa_1
Xfanout1412 fanout1419/X VGND VGND VPWR VPWR U$$2541/B sky130_fd_sc_hd__buf_8
Xfanout1423 U$$821/A VGND VGND VPWR VPWR U$$822/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1434 fanout1438/X VGND VGND VPWR VPWR U$$2412/B sky130_fd_sc_hd__buf_6
Xfanout1445 U$$2273/B VGND VGND VPWR VPWR U$$2301/B sky130_fd_sc_hd__buf_4
Xfanout1456 U$$2186/B VGND VGND VPWR VPWR U$$2191/A sky130_fd_sc_hd__buf_6
Xfanout1467 input22/X VGND VGND VPWR VPWR U$$2054/A sky130_fd_sc_hd__buf_6
XFILLER_65_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1041 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1478 U$$1727/B VGND VGND VPWR VPWR U$$1699/B sky130_fd_sc_hd__buf_4
Xfanout480 U$$3692/A2 VGND VGND VPWR VPWR U$$3696/A2 sky130_fd_sc_hd__buf_4
XFILLER_120_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1489 U$$1584/B VGND VGND VPWR VPWR U$$1570/B sky130_fd_sc_hd__buf_6
Xfanout491 U$$3439/A2 VGND VGND VPWR VPWR U$$3557/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_6_38_0 dadda_fa_6_38_0/A dadda_fa_6_38_0/B dadda_fa_6_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_39_0/B dadda_fa_7_38_0/CIN sky130_fd_sc_hd__fa_1
XU$$3203 U$$4162/A1 U$$3207/A2 U$$4162/B1 U$$3207/B2 VGND VGND VPWR VPWR U$$3204/A
+ sky130_fd_sc_hd__a22o_1
XU$$3214 U$$3214/A U$$3258/B VGND VGND VPWR VPWR U$$3214/X sky130_fd_sc_hd__xor2_1
XFILLER_171_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3225 U$$3499/A1 U$$3241/A2 U$$3636/B1 U$$3241/B2 VGND VGND VPWR VPWR U$$3226/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3236 U$$3236/A U$$3242/B VGND VGND VPWR VPWR U$$3236/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$18 _314_/Q _186_/Q VGND VGND VPWR VPWR final_adder.U$$237/A2 final_adder.U$$236/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3247 U$$3382/B1 U$$3251/A2 U$$3249/A1 U$$3251/B2 VGND VGND VPWR VPWR U$$3248/A
+ sky130_fd_sc_hd__a22o_1
XU$$2502 U$$447/A1 U$$2546/A2 U$$447/B1 U$$2546/B2 VGND VGND VPWR VPWR U$$2503/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$29 _325_/Q _197_/Q VGND VGND VPWR VPWR final_adder.U$$227/B1 final_adder.U$$226/B
+ sky130_fd_sc_hd__ha_1
XU$$3258 U$$3258/A U$$3258/B VGND VGND VPWR VPWR U$$3258/X sky130_fd_sc_hd__xor2_1
XU$$2513 U$$2513/A U$$2549/B VGND VGND VPWR VPWR U$$2513/X sky130_fd_sc_hd__xor2_1
XU$$2524 U$$3072/A1 U$$2532/A2 U$$3072/B1 U$$2532/B2 VGND VGND VPWR VPWR U$$2525/A
+ sky130_fd_sc_hd__a22o_1
XU$$3269 U$$3817/A1 U$$3285/A2 U$$3817/B1 U$$3285/B2 VGND VGND VPWR VPWR U$$3270/A
+ sky130_fd_sc_hd__a22o_1
XU$$2535 U$$2535/A U$$2541/B VGND VGND VPWR VPWR U$$2535/X sky130_fd_sc_hd__xor2_1
XU$$1801 U$$840/B1 U$$1841/A2 U$$707/A1 U$$1841/B2 VGND VGND VPWR VPWR U$$1802/A sky130_fd_sc_hd__a22o_1
XU$$2546 U$$80/A1 U$$2546/A2 U$$80/B1 U$$2546/B2 VGND VGND VPWR VPWR U$$2547/A sky130_fd_sc_hd__a22o_1
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2557 U$$2557/A U$$2603/A VGND VGND VPWR VPWR U$$2557/X sky130_fd_sc_hd__xor2_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1812 U$$1812/A U$$1836/B VGND VGND VPWR VPWR U$$1812/X sky130_fd_sc_hd__xor2_1
XU$$2568 U$$2840/B1 U$$2574/A2 U$$2707/A1 U$$2574/B2 VGND VGND VPWR VPWR U$$2569/A
+ sky130_fd_sc_hd__a22o_1
XU$$1823 U$$864/A1 U$$1829/A2 U$$864/B1 U$$1829/B2 VGND VGND VPWR VPWR U$$1824/A sky130_fd_sc_hd__a22o_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1834 U$$1834/A U$$1836/B VGND VGND VPWR VPWR U$$1834/X sky130_fd_sc_hd__xor2_1
XU$$2579 U$$2579/A U$$2603/A VGND VGND VPWR VPWR U$$2579/X sky130_fd_sc_hd__xor2_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1845 U$$612/A1 U$$1881/A2 U$$612/B1 U$$1881/B2 VGND VGND VPWR VPWR U$$1846/A sky130_fd_sc_hd__a22o_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1856 U$$1856/A U$$1882/B VGND VGND VPWR VPWR U$$1856/X sky130_fd_sc_hd__xor2_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1867 U$$3509/B1 U$$1909/A2 U$$3376/A1 U$$1909/B2 VGND VGND VPWR VPWR U$$1868/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1878 U$$1878/A U$$1916/B VGND VGND VPWR VPWR U$$1878/X sky130_fd_sc_hd__xor2_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1889 U$$654/B1 U$$1891/A2 U$$521/A1 U$$1891/B2 VGND VGND VPWR VPWR U$$1890/A sky130_fd_sc_hd__a22o_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_329_ _344_/CLK _329_/D VGND VGND VPWR VPWR _329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_70_2 dadda_fa_2_70_2/A dadda_fa_2_70_2/B dadda_fa_2_70_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_1/A dadda_fa_3_70_3/A sky130_fd_sc_hd__fa_1
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_63_1 dadda_fa_2_63_1/A dadda_fa_2_63_1/B dadda_fa_2_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_0/CIN dadda_fa_3_63_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$508 final_adder.U$$516/B final_adder.U$$508/B VGND VGND VPWR VPWR
+ final_adder.U$$628/B sky130_fd_sc_hd__and2_1
XFILLER_29_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$519 final_adder.U$$518/B final_adder.U$$403/X final_adder.U$$395/X
+ VGND VGND VPWR VPWR final_adder.U$$519/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_5_40_0 dadda_fa_5_40_0/A dadda_fa_5_40_0/B dadda_fa_5_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_41_0/A dadda_fa_6_40_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_56_0 dadda_fa_2_56_0/A dadda_fa_2_56_0/B dadda_fa_2_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_0/B dadda_fa_3_56_2/B sky130_fd_sc_hd__fa_1
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4460 U$$4460/A1 U$$4388/X U$$4460/B1 U$$4488/B2 VGND VGND VPWR VPWR U$$4461/A
+ sky130_fd_sc_hd__a22o_1
XU$$4471 U$$4471/A U$$4471/B VGND VGND VPWR VPWR U$$4471/X sky130_fd_sc_hd__xor2_1
XFILLER_53_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4482 U$$4482/A1 U$$4388/X U$$4482/B1 U$$4506/B2 VGND VGND VPWR VPWR U$$4483/A
+ sky130_fd_sc_hd__a22o_1
XU$$4493 U$$4493/A U$$4493/B VGND VGND VPWR VPWR U$$4493/X sky130_fd_sc_hd__xor2_1
XU$$3770 U$$3770/A U$$3774/B VGND VGND VPWR VPWR U$$3770/X sky130_fd_sc_hd__xor2_1
XU$$3781 U$$4466/A1 U$$3829/A2 U$$4468/A1 U$$3829/B2 VGND VGND VPWR VPWR U$$3782/A
+ sky130_fd_sc_hd__a22o_1
XU$$3792 U$$3792/A U$$3792/B VGND VGND VPWR VPWR U$$3792/X sky130_fd_sc_hd__xor2_1
XFILLER_40_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_85_2 dadda_fa_4_85_2/A dadda_fa_4_85_2/B dadda_fa_4_85_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_86_0/CIN dadda_fa_5_85_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_954 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_78_1 dadda_fa_4_78_1/A dadda_fa_4_78_1/B dadda_fa_4_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_79_0/B dadda_fa_5_78_1/B sky130_fd_sc_hd__fa_1
XFILLER_125_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_55_0 dadda_fa_7_55_0/A dadda_fa_7_55_0/B dadda_fa_7_55_0/CIN VGND VGND
+ VPWR VPWR _352_/D _223_/D sky130_fd_sc_hd__fa_1
XFILLER_115_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$903 U$$903/A U$$955/B VGND VGND VPWR VPWR U$$903/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_4_122_0_1946 VGND VGND VPWR VPWR dadda_ha_4_122_0/A dadda_ha_4_122_0_1946/LO
+ sky130_fd_sc_hd__conb_1
XU$$914 U$$914/A1 U$$956/A2 U$$914/B1 U$$956/B2 VGND VGND VPWR VPWR U$$915/A sky130_fd_sc_hd__a22o_1
XU$$925 U$$925/A U$$925/B VGND VGND VPWR VPWR U$$925/X sky130_fd_sc_hd__xor2_1
XFILLER_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$936 U$$936/A1 U$$942/A2 U$$936/B1 U$$942/B2 VGND VGND VPWR VPWR U$$937/A sky130_fd_sc_hd__a22o_1
XFILLER_84_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$947 U$$947/A U$$958/A VGND VGND VPWR VPWR U$$947/X sky130_fd_sc_hd__xor2_1
XU$$958 U$$958/A VGND VGND VPWR VPWR U$$958/Y sky130_fd_sc_hd__inv_1
XFILLER_43_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1108 U$$3298/B1 U$$1170/A2 U$$2480/A1 U$$1170/B2 VGND VGND VPWR VPWR U$$1109/A
+ sky130_fd_sc_hd__a22o_1
XU$$969 U$$969/A1 U$$981/A2 U$$971/A1 U$$981/B2 VGND VGND VPWR VPWR U$$970/A sky130_fd_sc_hd__a22o_1
XFILLER_55_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1119 U$$1119/A U$$1195/B VGND VGND VPWR VPWR U$$1119/X sky130_fd_sc_hd__xor2_1
XFILLER_141_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_80_1 dadda_fa_3_80_1/A dadda_fa_3_80_1/B dadda_fa_3_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_0/CIN dadda_fa_4_80_2/A sky130_fd_sc_hd__fa_1
XFILLER_152_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_73_0 dadda_fa_3_73_0/A dadda_fa_3_73_0/B dadda_fa_3_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_0/B dadda_fa_4_73_1/CIN sky130_fd_sc_hd__fa_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1220 U$$987/B1 VGND VGND VPWR VPWR U$$4001/B1 sky130_fd_sc_hd__buf_4
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1231 U$$3314/B1 VGND VGND VPWR VPWR U$$28/A1 sky130_fd_sc_hd__buf_4
Xfanout1242 input65/X VGND VGND VPWR VPWR U$$3979/B1 sky130_fd_sc_hd__buf_6
Xfanout1253 U$$547/A VGND VGND VPWR VPWR U$$504/B sky130_fd_sc_hd__buf_6
XFILLER_67_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1264 input60/X VGND VGND VPWR VPWR U$$4383/A sky130_fd_sc_hd__buf_4
XFILLER_66_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1275 fanout1279/X VGND VGND VPWR VPWR U$$4241/B sky130_fd_sc_hd__buf_2
Xfanout1286 U$$347/B VGND VGND VPWR VPWR U$$341/B sky130_fd_sc_hd__clkbuf_4
XU$$3000 U$$3000/A U$$3004/B VGND VGND VPWR VPWR U$$3000/X sky130_fd_sc_hd__xor2_1
Xfanout1297 U$$4058/B VGND VGND VPWR VPWR U$$4094/B sky130_fd_sc_hd__clkbuf_4
XU$$3011 U$$3285/A1 U$$3011/A2 U$$3011/B1 U$$3011/B2 VGND VGND VPWR VPWR U$$3012/A
+ sky130_fd_sc_hd__a22o_1
XU$$3022 U$$3022/A1 U$$3066/A2 U$$3022/B1 U$$3066/B2 VGND VGND VPWR VPWR U$$3023/A
+ sky130_fd_sc_hd__a22o_1
XU$$3033 U$$3033/A U$$3077/B VGND VGND VPWR VPWR U$$3033/X sky130_fd_sc_hd__xor2_1
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3044 U$$3181/A1 U$$3124/A2 U$$3181/B1 U$$3124/B2 VGND VGND VPWR VPWR U$$3045/A
+ sky130_fd_sc_hd__a22o_1
XU$$3055 U$$3055/A U$$3061/B VGND VGND VPWR VPWR U$$3055/X sky130_fd_sc_hd__xor2_1
XU$$2310 U$$2310/A1 U$$2310/A2 U$$2312/A1 U$$2310/B2 VGND VGND VPWR VPWR U$$2311/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_102_0 dadda_fa_4_102_0/A dadda_fa_4_102_0/B dadda_fa_4_102_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_103_0/A dadda_fa_5_102_1/A sky130_fd_sc_hd__fa_1
XU$$3066 U$$4162/A1 U$$3066/A2 U$$4162/B1 U$$3066/B2 VGND VGND VPWR VPWR U$$3067/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_35_5 U$$2338/X input185/X dadda_fa_2_35_5/CIN VGND VGND VPWR VPWR dadda_fa_3_36_2/A
+ dadda_fa_4_35_0/A sky130_fd_sc_hd__fa_2
XU$$2321 U$$2321/A U$$2327/B VGND VGND VPWR VPWR U$$2321/X sky130_fd_sc_hd__xor2_1
XU$$2332 U$$2446/B U$$2332/B VGND VGND VPWR VPWR U$$2332/X sky130_fd_sc_hd__and2_1
XU$$3077 U$$3077/A U$$3077/B VGND VGND VPWR VPWR U$$3077/X sky130_fd_sc_hd__xor2_1
XFILLER_34_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2343 U$$973/A1 U$$2415/A2 U$$973/B1 U$$2415/B2 VGND VGND VPWR VPWR U$$2344/A sky130_fd_sc_hd__a22o_1
XU$$3088 U$$4456/B1 U$$3112/A2 U$$4049/A1 U$$3112/B2 VGND VGND VPWR VPWR U$$3089/A
+ sky130_fd_sc_hd__a22o_1
XU$$2354 U$$2354/A U$$2396/B VGND VGND VPWR VPWR U$$2354/X sky130_fd_sc_hd__xor2_1
XU$$3099 U$$3099/A U$$3107/B VGND VGND VPWR VPWR U$$3099/X sky130_fd_sc_hd__xor2_1
XFILLER_62_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2365 U$$3322/B1 U$$2407/A2 U$$721/B1 U$$2407/B2 VGND VGND VPWR VPWR U$$2366/A
+ sky130_fd_sc_hd__a22o_1
XU$$1620 U$$1620/A U$$1626/B VGND VGND VPWR VPWR U$$1620/X sky130_fd_sc_hd__xor2_1
XU$$1631 U$$672/A1 U$$1641/A2 U$$672/B1 U$$1641/B2 VGND VGND VPWR VPWR U$$1632/A sky130_fd_sc_hd__a22o_1
XU$$2376 U$$2376/A U$$2416/B VGND VGND VPWR VPWR U$$2376/X sky130_fd_sc_hd__xor2_1
XU$$1642 U$$1642/A U$$1644/A VGND VGND VPWR VPWR U$$1642/X sky130_fd_sc_hd__xor2_1
XFILLER_50_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2387 U$$3072/A1 U$$2407/A2 U$$3072/B1 U$$2407/B2 VGND VGND VPWR VPWR U$$2388/A
+ sky130_fd_sc_hd__a22o_1
XU$$2398 U$$2398/A U$$2402/B VGND VGND VPWR VPWR U$$2398/X sky130_fd_sc_hd__xor2_1
XU$$1653 U$$1653/A U$$1699/B VGND VGND VPWR VPWR U$$1653/X sky130_fd_sc_hd__xor2_1
XU$$1664 U$$2897/A1 U$$1698/A2 U$$2897/B1 U$$1698/B2 VGND VGND VPWR VPWR U$$1665/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1675 U$$1675/A U$$1703/B VGND VGND VPWR VPWR U$$1675/X sky130_fd_sc_hd__xor2_1
XU$$1686 U$$864/A1 U$$1696/A2 U$$864/B1 U$$1696/B2 VGND VGND VPWR VPWR U$$1687/A sky130_fd_sc_hd__a22o_1
XU$$1697 U$$1697/A U$$1697/B VGND VGND VPWR VPWR U$$1697/X sky130_fd_sc_hd__xor2_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_95_1 dadda_fa_5_95_1/A dadda_fa_5_95_1/B dadda_fa_5_95_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_96_0/B dadda_fa_7_95_0/A sky130_fd_sc_hd__fa_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_88_0 dadda_fa_5_88_0/A dadda_fa_5_88_0/B dadda_fa_5_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_89_0/A dadda_fa_6_88_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_144_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$305 final_adder.U$$304/B final_adder.U$$179/X final_adder.U$$177/X
+ VGND VGND VPWR VPWR final_adder.U$$305/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$316 final_adder.U$$318/B final_adder.U$$316/B VGND VGND VPWR VPWR
+ final_adder.U$$442/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$327 final_adder.U$$326/B final_adder.U$$201/X final_adder.U$$199/X
+ VGND VGND VPWR VPWR final_adder.U$$327/X sky130_fd_sc_hd__a21o_1
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$338 final_adder.U$$340/B final_adder.U$$338/B VGND VGND VPWR VPWR
+ final_adder.U$$464/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$349 final_adder.U$$348/B final_adder.U$$223/X final_adder.U$$221/X
+ VGND VGND VPWR VPWR final_adder.U$$349/X sky130_fd_sc_hd__a21o_1
XFILLER_26_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4290 U$$4290/A U$$4383/A VGND VGND VPWR VPWR U$$4290/X sky130_fd_sc_hd__xor2_1
XFILLER_38_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4401_1848 VGND VGND VPWR VPWR U$$4401_1848/HI U$$4401/B sky130_fd_sc_hd__conb_1
Xdadda_fa_4_90_0 dadda_fa_4_90_0/A dadda_fa_4_90_0/B dadda_fa_4_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_91_0/A dadda_fa_5_90_1/A sky130_fd_sc_hd__fa_1
XFILLER_107_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_104_2 input134/X dadda_fa_3_104_2/B dadda_fa_3_104_2/CIN VGND VGND VPWR
+ VPWR dadda_fa_4_105_1/A dadda_fa_4_104_2/B sky130_fd_sc_hd__fa_1
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_118_0 dadda_fa_6_118_0/A dadda_fa_6_118_0/B dadda_fa_6_118_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_119_0/B dadda_fa_7_118_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$861 final_adder.U$$764/X final_adder.U$$829/X final_adder.U$$765/X
+ VGND VGND VPWR VPWR final_adder.U$$861/X sky130_fd_sc_hd__a21o_2
XU$$700 U$$700/A U$$744/B VGND VGND VPWR VPWR U$$700/X sky130_fd_sc_hd__xor2_1
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$711 U$$26/A1 U$$743/A2 U$$28/A1 U$$743/B2 VGND VGND VPWR VPWR U$$712/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$883 final_adder.U$$786/X final_adder.U$$619/X final_adder.U$$787/X
+ VGND VGND VPWR VPWR final_adder.U$$883/X sky130_fd_sc_hd__a21o_1
XU$$722 U$$722/A U$$768/B VGND VGND VPWR VPWR U$$722/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_38_3 dadda_fa_3_38_3/A dadda_fa_3_38_3/B dadda_fa_3_38_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_1/B dadda_fa_4_38_2/CIN sky130_fd_sc_hd__fa_1
XU$$733 U$$868/B1 U$$769/A2 U$$735/A1 U$$769/B2 VGND VGND VPWR VPWR U$$734/A sky130_fd_sc_hd__a22o_1
XFILLER_17_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$744 U$$744/A U$$744/B VGND VGND VPWR VPWR U$$744/X sky130_fd_sc_hd__xor2_1
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$755 U$$892/A1 U$$763/A2 U$$894/A1 U$$763/B2 VGND VGND VPWR VPWR U$$756/A sky130_fd_sc_hd__a22o_1
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$766 U$$766/A U$$768/B VGND VGND VPWR VPWR U$$766/X sky130_fd_sc_hd__xor2_1
XFILLER_72_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$777 U$$914/A1 U$$819/A2 U$$914/B1 U$$819/B2 VGND VGND VPWR VPWR U$$778/A sky130_fd_sc_hd__a22o_1
XU$$788 U$$788/A U$$820/B VGND VGND VPWR VPWR U$$788/X sky130_fd_sc_hd__xor2_1
XFILLER_31_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$799 U$$936/A1 U$$809/A2 U$$936/B1 U$$809/B2 VGND VGND VPWR VPWR U$$800/A sky130_fd_sc_hd__a22o_1
XFILLER_16_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1050 U$$3846/B1 VGND VGND VPWR VPWR U$$697/A1 sky130_fd_sc_hd__buf_2
XFILLER_6_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1061 input86/X VGND VGND VPWR VPWR U$$3080/A1 sky130_fd_sc_hd__buf_6
Xfanout1072 input84/X VGND VGND VPWR VPWR U$$2665/A1 sky130_fd_sc_hd__buf_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1083 U$$4442/B1 VGND VGND VPWR VPWR U$$4307/A1 sky130_fd_sc_hd__buf_4
Xfanout1094 U$$56/A1 VGND VGND VPWR VPWR U$$465/B1 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_2_40_3 U$$2747/X U$$2805/B input191/X VGND VGND VPWR VPWR dadda_fa_3_41_1/B
+ dadda_fa_3_40_3/B sky130_fd_sc_hd__fa_1
XFILLER_19_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_33_2 U$$871/X U$$1004/X U$$1137/X VGND VGND VPWR VPWR dadda_fa_3_34_1/A
+ dadda_fa_3_33_3/A sky130_fd_sc_hd__fa_1
XU$$2140 U$$2140/A U$$2140/B VGND VGND VPWR VPWR U$$2140/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_10_1 dadda_fa_5_10_1/A dadda_fa_5_10_1/B dadda_ha_4_10_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_11_0/B dadda_fa_7_10_0/A sky130_fd_sc_hd__fa_1
XU$$2151 U$$3382/B1 U$$2189/A2 U$$3249/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2152/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_26_1 U$$458/X U$$591/X U$$724/X VGND VGND VPWR VPWR dadda_fa_3_27_2/CIN
+ dadda_fa_3_26_3/CIN sky130_fd_sc_hd__fa_1
XU$$2162 U$$2162/A U$$2192/A VGND VGND VPWR VPWR U$$2162/X sky130_fd_sc_hd__xor2_1
XU$$2173 U$$2310/A1 U$$2181/A2 U$$2312/A1 U$$2181/B2 VGND VGND VPWR VPWR U$$2174/A
+ sky130_fd_sc_hd__a22o_1
XU$$2184 U$$2184/A U$$2186/B VGND VGND VPWR VPWR U$$2184/X sky130_fd_sc_hd__xor2_1
XU$$2195 U$$2329/A U$$2195/B VGND VGND VPWR VPWR U$$2195/X sky130_fd_sc_hd__and2_1
XU$$1450 U$$80/A1 U$$1452/A2 U$$80/B1 U$$1452/B2 VGND VGND VPWR VPWR U$$1451/A sky130_fd_sc_hd__a22o_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1461 U$$1461/A U$$1461/B VGND VGND VPWR VPWR U$$1461/X sky130_fd_sc_hd__xor2_1
XU$$1472 U$$924/A1 U$$1504/A2 U$$2979/B1 U$$1504/B2 VGND VGND VPWR VPWR U$$1473/A
+ sky130_fd_sc_hd__a22o_1
XU$$1483 U$$1483/A U$$1491/B VGND VGND VPWR VPWR U$$1483/X sky130_fd_sc_hd__xor2_1
XFILLER_148_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1494 U$$2042/A1 U$$1504/A2 U$$2179/B1 U$$1504/B2 VGND VGND VPWR VPWR U$$1495/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_85_5 U$$3502/X U$$3635/X U$$3768/X VGND VGND VPWR VPWR dadda_fa_2_86_4/A
+ dadda_fa_3_85_0/A sky130_fd_sc_hd__fa_2
XFILLER_132_957 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_78_4 U$$2823/X U$$2956/X U$$3089/X VGND VGND VPWR VPWR dadda_fa_2_79_1/CIN
+ dadda_fa_2_78_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_170_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$102 _398_/Q _270_/Q VGND VGND VPWR VPWR final_adder.U$$923/B1 final_adder.U$$152/A
+ sky130_fd_sc_hd__ha_1
XFILLER_100_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$113 _409_/Q _281_/Q VGND VGND VPWR VPWR final_adder.U$$143/B1 final_adder.U$$142/B
+ sky130_fd_sc_hd__ha_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_48_2 dadda_fa_4_48_2/A dadda_fa_4_48_2/B dadda_fa_4_48_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_49_0/CIN dadda_fa_5_48_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$124 _420_/Q _292_/Q VGND VGND VPWR VPWR final_adder.U$$901/B1 final_adder.U$$130/A
+ sky130_fd_sc_hd__ha_1
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$135 final_adder.U$$134/B final_adder.U$$905/B1 final_adder.U$$135/B1
+ VGND VGND VPWR VPWR final_adder.U$$135/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$146 final_adder.U$$146/A final_adder.U$$146/B VGND VGND VPWR VPWR
+ final_adder.U$$274/B sky130_fd_sc_hd__and2_1
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$157 final_adder.U$$156/B final_adder.U$$927/B1 final_adder.U$$157/B1
+ VGND VGND VPWR VPWR final_adder.U$$157/X sky130_fd_sc_hd__a21o_1
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$168 final_adder.U$$168/A final_adder.U$$168/B VGND VGND VPWR VPWR
+ final_adder.U$$296/B sky130_fd_sc_hd__and2_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$179 final_adder.U$$178/B final_adder.U$$949/B1 final_adder.U$$179/B1
+ VGND VGND VPWR VPWR final_adder.U$$179/X sky130_fd_sc_hd__a21o_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_18_0 dadda_fa_7_18_0/A dadda_fa_7_18_0/B dadda_fa_7_18_0/CIN VGND VGND
+ VPWR VPWR _315_/D _186_/D sky130_fd_sc_hd__fa_2
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4399_1847 VGND VGND VPWR VPWR U$$4399_1847/HI U$$4399/B sky130_fd_sc_hd__conb_1
XFILLER_127_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput120 b[5] VGND VGND VPWR VPWR input120/X sky130_fd_sc_hd__buf_4
Xinput131 c[101] VGND VGND VPWR VPWR input131/X sky130_fd_sc_hd__buf_4
XFILLER_0_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_50_2 dadda_fa_3_50_2/A dadda_fa_3_50_2/B dadda_fa_3_50_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_1/A dadda_fa_4_50_2/B sky130_fd_sc_hd__fa_1
XFILLER_103_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput142 c[111] VGND VGND VPWR VPWR input142/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_0_66_2 U$$937/X U$$1070/X U$$1203/X VGND VGND VPWR VPWR dadda_fa_1_67_6/A
+ dadda_fa_1_66_8/A sky130_fd_sc_hd__fa_1
Xinput153 c[121] VGND VGND VPWR VPWR input153/X sky130_fd_sc_hd__buf_2
Xinput164 c[16] VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__buf_2
Xinput175 c[26] VGND VGND VPWR VPWR input175/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_3_43_1 dadda_fa_3_43_1/A dadda_fa_3_43_1/B dadda_fa_3_43_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_0/CIN dadda_fa_4_43_2/A sky130_fd_sc_hd__fa_1
Xinput186 c[36] VGND VGND VPWR VPWR input186/X sky130_fd_sc_hd__clkbuf_4
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_59_1 U$$524/X U$$657/X U$$790/X VGND VGND VPWR VPWR dadda_fa_1_60_6/CIN
+ dadda_fa_1_59_8/B sky130_fd_sc_hd__fa_2
XFILLER_56_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput197 c[46] VGND VGND VPWR VPWR input197/X sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_6_20_0 dadda_fa_6_20_0/A dadda_fa_6_20_0/B dadda_fa_6_20_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_21_0/B dadda_fa_7_20_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$680 final_adder.U$$696/B final_adder.U$$680/B VGND VGND VPWR VPWR
+ final_adder.U$$792/B sky130_fd_sc_hd__and2_1
Xdadda_fa_3_36_0 dadda_fa_3_36_0/A dadda_fa_3_36_0/B dadda_fa_3_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_0/B dadda_fa_4_36_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$691 final_adder.U$$690/B final_adder.U$$587/X final_adder.U$$571/X
+ VGND VGND VPWR VPWR final_adder.U$$691/X sky130_fd_sc_hd__a21o_1
XU$$530 U$$530/A U$$536/B VGND VGND VPWR VPWR U$$530/X sky130_fd_sc_hd__xor2_1
XU$$541 U$$678/A1 U$$543/A2 U$$678/B1 U$$543/B2 VGND VGND VPWR VPWR U$$542/A sky130_fd_sc_hd__a22o_1
XU$$552 U$$550/Y U$$549/A U$$548/A U$$551/X U$$548/Y VGND VGND VPWR VPWR U$$552/X
+ sky130_fd_sc_hd__a32o_2
XU$$563 U$$563/A U$$643/B VGND VGND VPWR VPWR U$$563/X sky130_fd_sc_hd__xor2_1
XFILLER_44_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$574 U$$709/B1 U$$638/A2 U$$576/A1 U$$638/B2 VGND VGND VPWR VPWR U$$575/A sky130_fd_sc_hd__a22o_1
XU$$585 U$$585/A U$$637/B VGND VGND VPWR VPWR U$$585/X sky130_fd_sc_hd__xor2_1
XU$$596 U$$596/A1 U$$630/A2 U$$596/B1 U$$630/B2 VGND VGND VPWR VPWR U$$597/A sky130_fd_sc_hd__a22o_1
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_95_4 U$$4187/X U$$4320/X U$$4453/X VGND VGND VPWR VPWR dadda_fa_3_96_1/CIN
+ dadda_fa_3_95_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_88_3 dadda_fa_2_88_3/A dadda_fa_2_88_3/B dadda_fa_2_88_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_89_1/B dadda_fa_3_88_3/B sky130_fd_sc_hd__fa_1
XFILLER_99_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_58_1 dadda_fa_5_58_1/A dadda_fa_5_58_1/B dadda_fa_5_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_59_0/B dadda_fa_7_58_0/A sky130_fd_sc_hd__fa_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_104_1 U$$3141/X U$$3274/X U$$3407/X VGND VGND VPWR VPWR dadda_fa_3_105_3/A
+ dadda_fa_3_104_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1280 U$$1280/A U$$1282/B VGND VGND VPWR VPWR U$$1280/X sky130_fd_sc_hd__xor2_1
XU$$1291 U$$58/A1 U$$1295/A2 U$$60/A1 U$$1295/B2 VGND VGND VPWR VPWR U$$1292/A sky130_fd_sc_hd__a22o_1
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_125_0 U$$4246/Y U$$4380/X U$$4513/X VGND VGND VPWR VPWR dadda_fa_6_126_0/CIN
+ dadda_fa_7_125_0/A sky130_fd_sc_hd__fa_1
XFILLER_164_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_2 U$$2168/X U$$2301/X U$$2434/X VGND VGND VPWR VPWR dadda_fa_2_84_2/B
+ dadda_fa_2_83_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_131_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout810 U$$2679/B2 VGND VGND VPWR VPWR U$$2733/B2 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_4_60_1 dadda_fa_4_60_1/A dadda_fa_4_60_1/B dadda_fa_4_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_61_0/B dadda_fa_5_60_1/B sky130_fd_sc_hd__fa_1
Xfanout821 U$$2407/B2 VGND VGND VPWR VPWR U$$2395/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_76_1 U$$1888/X U$$2021/X U$$2154/X VGND VGND VPWR VPWR dadda_fa_2_77_0/CIN
+ dadda_fa_2_76_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout832 U$$2282/B2 VGND VGND VPWR VPWR U$$2248/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout843 U$$2060/X VGND VGND VPWR VPWR U$$2181/B2 sky130_fd_sc_hd__buf_6
Xfanout854 U$$1859/B2 VGND VGND VPWR VPWR U$$1831/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_53_0 dadda_fa_4_53_0/A dadda_fa_4_53_0/B dadda_fa_4_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_54_0/A dadda_fa_5_53_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_69_0 U$$2406/X U$$2539/X U$$2672/X VGND VGND VPWR VPWR dadda_fa_2_70_0/B
+ dadda_fa_2_69_3/B sky130_fd_sc_hd__fa_1
Xfanout865 U$$1720/B2 VGND VGND VPWR VPWR U$$1702/B2 sky130_fd_sc_hd__buf_4
Xfanout876 U$$1625/B2 VGND VGND VPWR VPWR U$$1641/B2 sky130_fd_sc_hd__clkbuf_8
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout887 U$$142/X VGND VGND VPWR VPWR U$$253/B2 sky130_fd_sc_hd__buf_6
Xfanout898 U$$1361/B2 VGND VGND VPWR VPWR U$$1367/B2 sky130_fd_sc_hd__buf_4
XFILLER_46_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2909 U$$4416/A1 U$$2989/A2 U$$4416/B1 U$$2989/B2 VGND VGND VPWR VPWR U$$2910/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_362_ _364_/CLK _362_/D VGND VGND VPWR VPWR _362_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_293_ _421_/CLK _293_/D VGND VGND VPWR VPWR _293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_98_2 dadda_fa_3_98_2/A dadda_fa_3_98_2/B dadda_fa_3_98_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_99_1/A dadda_fa_4_98_2/B sky130_fd_sc_hd__fa_1
XFILLER_107_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_68_0 dadda_fa_6_68_0/A dadda_fa_6_68_0/B dadda_fa_6_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_69_0/B dadda_fa_7_68_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_123_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4453_1874 VGND VGND VPWR VPWR U$$4453_1874/HI U$$4453/B sky130_fd_sc_hd__conb_1
XFILLER_111_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_71_0 U$$547/Y U$$681/X U$$814/X VGND VGND VPWR VPWR dadda_fa_1_72_6/CIN
+ dadda_fa_1_71_8/A sky130_fd_sc_hd__fa_1
XFILLER_49_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_5_7_1 U$$420/X input234/X VGND VGND VPWR VPWR dadda_fa_6_8_0/B dadda_fa_7_7_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_91_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$360 U$$632/B1 U$$362/A2 U$$499/A1 U$$362/B2 VGND VGND VPWR VPWR U$$361/A sky130_fd_sc_hd__a22o_1
XFILLER_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$371 U$$371/A U$$410/A VGND VGND VPWR VPWR U$$371/X sky130_fd_sc_hd__xor2_1
XU$$382 U$$517/B1 U$$386/A2 U$$384/A1 U$$386/B2 VGND VGND VPWR VPWR U$$383/A sky130_fd_sc_hd__a22o_1
XU$$393 U$$393/A U$$410/A VGND VGND VPWR VPWR U$$393/X sky130_fd_sc_hd__xor2_1
XFILLER_33_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_93_1 U$$3252/X U$$3385/X U$$3518/X VGND VGND VPWR VPWR dadda_fa_3_94_0/CIN
+ dadda_fa_3_93_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_70_0 dadda_fa_5_70_0/A dadda_fa_5_70_0/B dadda_fa_5_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_71_0/A dadda_fa_6_70_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_86_0 U$$3770/X U$$3903/X U$$4036/X VGND VGND VPWR VPWR dadda_fa_3_87_0/B
+ dadda_fa_3_86_2/B sky130_fd_sc_hd__fa_1
XFILLER_141_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_49_7 U$$2898/X U$$3031/X VGND VGND VPWR VPWR dadda_fa_2_50_3/A dadda_fa_3_49_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_87_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_62_7 dadda_fa_1_62_7/A dadda_fa_1_62_7/B dadda_fa_1_62_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_63_2/CIN dadda_fa_2_62_5/CIN sky130_fd_sc_hd__fa_1
XU$$1924_1796 VGND VGND VPWR VPWR U$$1924_1796/HI U$$1924/A1 sky130_fd_sc_hd__conb_1
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_55_6 U$$3176/X U$$3309/X U$$3442/X VGND VGND VPWR VPWR dadda_fa_2_56_2/B
+ dadda_fa_2_55_5/B sky130_fd_sc_hd__fa_1
XFILLER_55_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_48_5 U$$2098/X U$$2231/X U$$2364/X VGND VGND VPWR VPWR dadda_fa_2_49_2/CIN
+ dadda_fa_2_48_5/B sky130_fd_sc_hd__fa_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_7_0 dadda_fa_7_7_0/A dadda_fa_7_7_0/B dadda_fa_7_7_0/CIN VGND VGND VPWR
+ VPWR _304_/D _175_/D sky130_fd_sc_hd__fa_1
XFILLER_36_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_944 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_85_0 dadda_fa_7_85_0/A dadda_fa_7_85_0/B dadda_fa_7_85_0/CIN VGND VGND
+ VPWR VPWR _382_/D _253_/D sky130_fd_sc_hd__fa_2
XFILLER_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1605 U$$4508/A1 VGND VGND VPWR VPWR U$$4234/A1 sky130_fd_sc_hd__buf_4
Xfanout1616 U$$4506/A1 VGND VGND VPWR VPWR U$$4093/B1 sky130_fd_sc_hd__buf_2
Xfanout1627 input116/X VGND VGND VPWR VPWR U$$2860/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout640 U$$1237/X VGND VGND VPWR VPWR U$$1361/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1638 U$$938/A1 VGND VGND VPWR VPWR U$$2443/B1 sky130_fd_sc_hd__buf_4
Xfanout1649 U$$2578/B1 VGND VGND VPWR VPWR U$$251/A1 sky130_fd_sc_hd__buf_2
Xfanout651 U$$1202/A2 VGND VGND VPWR VPWR U$$1218/A2 sky130_fd_sc_hd__buf_6
Xfanout662 U$$952/B2 VGND VGND VPWR VPWR U$$942/B2 sky130_fd_sc_hd__buf_6
XU$$4108 U$$4108/A U$$4108/B VGND VGND VPWR VPWR U$$4108/X sky130_fd_sc_hd__xor2_1
XU$$4119 U$$4119/A U$$4133/B VGND VGND VPWR VPWR U$$4119/X sky130_fd_sc_hd__xor2_1
Xfanout673 U$$819/B2 VGND VGND VPWR VPWR U$$771/B2 sky130_fd_sc_hd__buf_4
Xfanout684 U$$4289/B2 VGND VGND VPWR VPWR U$$4295/B2 sky130_fd_sc_hd__buf_4
Xfanout695 U$$543/B2 VGND VGND VPWR VPWR U$$539/B2 sky130_fd_sc_hd__buf_4
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3407 U$$3407/A U$$3411/B VGND VGND VPWR VPWR U$$3407/X sky130_fd_sc_hd__xor2_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3418 U$$3418/A1 U$$3418/A2 U$$3418/B1 U$$3418/B2 VGND VGND VPWR VPWR U$$3419/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_100_0 dadda_fa_6_100_0/A dadda_fa_6_100_0/B dadda_fa_6_100_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_101_0/B dadda_fa_7_100_0/CIN sky130_fd_sc_hd__fa_1
XU$$3429 U$$3427/Y input46/X U$$3425/A U$$3428/X U$$3425/Y VGND VGND VPWR VPWR U$$3429/X
+ sky130_fd_sc_hd__a32o_2
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2706 U$$2706/A U$$2708/B VGND VGND VPWR VPWR U$$2706/X sky130_fd_sc_hd__xor2_1
XFILLER_46_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2717 U$$4361/A1 U$$2733/A2 U$$4363/A1 U$$2733/B2 VGND VGND VPWR VPWR U$$2718/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2728 U$$2728/A U$$2738/B VGND VGND VPWR VPWR U$$2728/X sky130_fd_sc_hd__xor2_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2739 U$$2739/A VGND VGND VPWR VPWR U$$2739/Y sky130_fd_sc_hd__inv_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4483_1889 VGND VGND VPWR VPWR U$$4483_1889/HI U$$4483/B sky130_fd_sc_hd__conb_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_414_ _421_/CLK _414_/D VGND VGND VPWR VPWR _414_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_345_ _345_/CLK _345_/D VGND VGND VPWR VPWR _345_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_276_ _405_/CLK _276_/D VGND VGND VPWR VPWR _276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_65_5 dadda_fa_2_65_5/A dadda_fa_2_65_5/B dadda_fa_2_65_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_2/A dadda_fa_4_65_0/A sky130_fd_sc_hd__fa_2
XFILLER_96_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_58_4 dadda_fa_2_58_4/A dadda_fa_2_58_4/B dadda_fa_2_58_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_1/CIN dadda_fa_3_58_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_110_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3930 U$$4341/A1 U$$3960/A2 U$$4480/A1 U$$3960/B2 VGND VGND VPWR VPWR U$$3931/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3941 U$$3941/A U$$3961/B VGND VGND VPWR VPWR U$$3941/X sky130_fd_sc_hd__xor2_1
XU$$3952 U$$4363/A1 U$$3966/A2 U$$4365/A1 U$$3966/B2 VGND VGND VPWR VPWR U$$3953/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3963 U$$3963/A U$$3965/B VGND VGND VPWR VPWR U$$3963/X sky130_fd_sc_hd__xor2_1
XU$$3974 input54/X VGND VGND VPWR VPWR U$$3976/B sky130_fd_sc_hd__inv_1
XFILLER_91_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3985 U$$4257/B1 U$$4025/A2 U$$4259/B1 U$$4025/B2 VGND VGND VPWR VPWR U$$3986/A
+ sky130_fd_sc_hd__a22o_1
XU$$3996 U$$3996/A U$$4026/B VGND VGND VPWR VPWR U$$3996/X sky130_fd_sc_hd__xor2_1
XFILLER_18_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$190 U$$190/A U$$220/B VGND VGND VPWR VPWR U$$190/X sky130_fd_sc_hd__xor2_1
XFILLER_33_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput265 output265/A VGND VGND VPWR VPWR o[107] sky130_fd_sc_hd__buf_2
Xoutput276 output276/A VGND VGND VPWR VPWR o[117] sky130_fd_sc_hd__buf_2
XFILLER_88_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput287 output287/A VGND VGND VPWR VPWR o[127] sky130_fd_sc_hd__buf_2
XFILLER_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput298 output298/A VGND VGND VPWR VPWR o[21] sky130_fd_sc_hd__buf_2
XFILLER_102_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_60_4 U$$3585/X U$$3718/X U$$3851/X VGND VGND VPWR VPWR dadda_fa_2_61_1/CIN
+ dadda_fa_2_60_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_3 U$$1576/X U$$1709/X U$$1842/X VGND VGND VPWR VPWR dadda_fa_2_54_1/B
+ dadda_fa_2_53_4/B sky130_fd_sc_hd__fa_1
XFILLER_56_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_30_2 dadda_fa_4_30_2/A dadda_fa_4_30_2/B dadda_fa_4_30_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_31_0/CIN dadda_fa_5_30_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_46_2 U$$897/X U$$1030/X U$$1163/X VGND VGND VPWR VPWR dadda_fa_2_47_2/B
+ dadda_fa_2_46_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_23_1 dadda_fa_4_23_1/A dadda_fa_4_23_1/B dadda_fa_4_23_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_24_0/B dadda_fa_5_23_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_39_1 U$$484/X U$$617/X U$$750/X VGND VGND VPWR VPWR dadda_fa_2_40_4/B
+ dadda_fa_2_39_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_167_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_16_0 U$$704/X U$$837/X U$$970/X VGND VGND VPWR VPWR dadda_fa_5_17_0/A
+ dadda_fa_5_16_1/A sky130_fd_sc_hd__fa_1
XFILLER_168_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1106 final_adder.U$$172/A final_adder.U$$881/X VGND VGND VPWR VPWR
+ output365/A sky130_fd_sc_hd__xor2_1
XFILLER_11_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1117 final_adder.U$$162/B final_adder.U$$933/X VGND VGND VPWR VPWR
+ output377/A sky130_fd_sc_hd__xor2_1
XFILLER_128_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1128 final_adder.U$$150/A final_adder.U$$859/X VGND VGND VPWR VPWR
+ output262/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1139 final_adder.U$$140/B final_adder.U$$911/X VGND VGND VPWR VPWR
+ output274/A sky130_fd_sc_hd__xor2_1
XFILLER_124_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1402 U$$2668/B VGND VGND VPWR VPWR U$$2662/B sky130_fd_sc_hd__buf_6
XFILLER_120_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1413 fanout1419/X VGND VGND VPWR VPWR U$$2575/B sky130_fd_sc_hd__buf_6
Xdadda_fa_3_68_3 dadda_fa_3_68_3/A dadda_fa_3_68_3/B dadda_fa_3_68_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_1/B dadda_fa_4_68_2/CIN sky130_fd_sc_hd__fa_1
Xfanout1424 U$$778/B VGND VGND VPWR VPWR U$$744/B sky130_fd_sc_hd__clkbuf_8
Xfanout1435 fanout1438/X VGND VGND VPWR VPWR U$$2416/B sky130_fd_sc_hd__buf_6
Xfanout1446 U$$2328/A VGND VGND VPWR VPWR U$$2327/B sky130_fd_sc_hd__buf_6
Xfanout1457 input25/X VGND VGND VPWR VPWR U$$2186/B sky130_fd_sc_hd__buf_4
Xfanout1468 U$$1832/B VGND VGND VPWR VPWR U$$1828/B sky130_fd_sc_hd__buf_6
Xfanout470 U$$3777/A2 VGND VGND VPWR VPWR U$$3773/A2 sky130_fd_sc_hd__buf_4
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout481 U$$3692/A2 VGND VGND VPWR VPWR U$$3682/A2 sky130_fd_sc_hd__buf_4
XFILLER_24_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1479 input18/X VGND VGND VPWR VPWR U$$1727/B sky130_fd_sc_hd__clkbuf_4
Xfanout492 U$$3429/X VGND VGND VPWR VPWR U$$3439/A2 sky130_fd_sc_hd__buf_6
XFILLER_59_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3204 U$$3204/A U$$3208/B VGND VGND VPWR VPWR U$$3204/X sky130_fd_sc_hd__xor2_1
XFILLER_46_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3215 U$$4446/B1 U$$3283/A2 U$$4450/A1 U$$3283/B2 VGND VGND VPWR VPWR U$$3216/A
+ sky130_fd_sc_hd__a22o_1
XU$$3226 U$$3226/A U$$3242/B VGND VGND VPWR VPWR U$$3226/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$19 _315_/Q _187_/Q VGND VGND VPWR VPWR final_adder.U$$237/B1 final_adder.U$$236/B
+ sky130_fd_sc_hd__ha_1
XFILLER_19_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3237 U$$3372/B1 U$$3241/A2 U$$3239/A1 U$$3241/B2 VGND VGND VPWR VPWR U$$3238/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3248 U$$3248/A U$$3287/A VGND VGND VPWR VPWR U$$3248/X sky130_fd_sc_hd__xor2_1
XU$$2503 U$$2503/A U$$2545/B VGND VGND VPWR VPWR U$$2503/X sky130_fd_sc_hd__xor2_1
XU$$3259 U$$4081/A1 U$$3283/A2 U$$4081/B1 U$$3283/B2 VGND VGND VPWR VPWR U$$3260/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2514 U$$870/A1 U$$2546/A2 U$$872/A1 U$$2546/B2 VGND VGND VPWR VPWR U$$2515/A sky130_fd_sc_hd__a22o_1
XU$$2525 U$$2525/A U$$2529/B VGND VGND VPWR VPWR U$$2525/X sky130_fd_sc_hd__xor2_1
XFILLER_73_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2536 U$$3630/B1 U$$2578/A2 U$$3495/B1 U$$2578/B2 VGND VGND VPWR VPWR U$$2537/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1802 U$$1802/A U$$1836/B VGND VGND VPWR VPWR U$$1802/X sky130_fd_sc_hd__xor2_1
XU$$2547 U$$2547/A U$$2549/B VGND VGND VPWR VPWR U$$2547/X sky130_fd_sc_hd__xor2_1
XU$$1813 U$$852/B1 U$$1841/A2 U$$34/A1 U$$1841/B2 VGND VGND VPWR VPWR U$$1814/A sky130_fd_sc_hd__a22o_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2558 U$$3243/A1 U$$2578/A2 U$$3243/B1 U$$2578/B2 VGND VGND VPWR VPWR U$$2559/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2569 U$$2569/A U$$2575/B VGND VGND VPWR VPWR U$$2569/X sky130_fd_sc_hd__xor2_1
XU$$1824 U$$1824/A U$$1828/B VGND VGND VPWR VPWR U$$1824/X sky130_fd_sc_hd__xor2_1
XFILLER_62_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1835 U$$739/A1 U$$1841/A2 U$$741/A1 U$$1841/B2 VGND VGND VPWR VPWR U$$1836/A sky130_fd_sc_hd__a22o_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1846 U$$1846/A U$$1854/B VGND VGND VPWR VPWR U$$1846/X sky130_fd_sc_hd__xor2_1
XU$$1857 U$$487/A1 U$$1859/A2 U$$487/B1 U$$1859/B2 VGND VGND VPWR VPWR U$$1858/A sky130_fd_sc_hd__a22o_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1868 U$$1868/A U$$1874/B VGND VGND VPWR VPWR U$$1868/X sky130_fd_sc_hd__xor2_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1879 U$$920/A1 U$$1915/A2 U$$920/B1 U$$1915/B2 VGND VGND VPWR VPWR U$$1880/A sky130_fd_sc_hd__a22o_1
XFILLER_159_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_328_ _328_/CLK _328_/D VGND VGND VPWR VPWR _328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_259_ _423_/CLK _259_/D VGND VGND VPWR VPWR _259_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_952 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_70_3 dadda_fa_2_70_3/A dadda_fa_2_70_3/B dadda_fa_2_70_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_1/B dadda_fa_3_70_3/B sky130_fd_sc_hd__fa_1
XFILLER_130_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_63_2 dadda_fa_2_63_2/A dadda_fa_2_63_2/B dadda_fa_2_63_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_1/A dadda_fa_3_63_3/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$509 final_adder.U$$508/B final_adder.U$$393/X final_adder.U$$385/X
+ VGND VGND VPWR VPWR final_adder.U$$509/X sky130_fd_sc_hd__a21o_1
XFILLER_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_40_1 dadda_fa_5_40_1/A dadda_fa_5_40_1/B dadda_fa_5_40_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_41_0/B dadda_fa_7_40_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_56_1 dadda_fa_2_56_1/A dadda_fa_2_56_1/B dadda_fa_2_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_0/CIN dadda_fa_3_56_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_33_0 dadda_fa_5_33_0/A dadda_fa_5_33_0/B dadda_fa_5_33_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_34_0/A dadda_fa_6_33_0/CIN sky130_fd_sc_hd__fa_2
XU$$4450 U$$4450/A1 U$$4388/X U$$4452/A1 U$$4458/B2 VGND VGND VPWR VPWR U$$4451/A
+ sky130_fd_sc_hd__a22o_1
XU$$4386_1838 VGND VGND VPWR VPWR U$$4386_1838/HI U$$4386/A sky130_fd_sc_hd__conb_1
XFILLER_49_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_49_0 U$$3164/X U$$3297/X input200/X VGND VGND VPWR VPWR dadda_fa_3_50_0/B
+ dadda_fa_3_49_2/B sky130_fd_sc_hd__fa_1
XU$$4461 U$$4461/A U$$4461/B VGND VGND VPWR VPWR U$$4461/X sky130_fd_sc_hd__xor2_1
XU$$4472 U$$4472/A1 U$$4388/X U$$4474/A1 U$$4492/B2 VGND VGND VPWR VPWR U$$4473/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4483 U$$4483/A U$$4483/B VGND VGND VPWR VPWR U$$4483/X sky130_fd_sc_hd__xor2_1
XFILLER_53_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4494 U$$4494/A1 U$$4388/X U$$4496/A1 U$$4506/B2 VGND VGND VPWR VPWR U$$4495/A
+ sky130_fd_sc_hd__a22o_1
XU$$3760 U$$3760/A U$$3774/B VGND VGND VPWR VPWR U$$3760/X sky130_fd_sc_hd__xor2_1
XU$$3771 U$$4043/B1 U$$3773/A2 U$$3908/B1 U$$3773/B2 VGND VGND VPWR VPWR U$$3772/A
+ sky130_fd_sc_hd__a22o_1
XU$$3782 U$$3782/A U$$3828/B VGND VGND VPWR VPWR U$$3782/X sky130_fd_sc_hd__xor2_1
XU$$3793 U$$4478/A1 U$$3825/A2 U$$4478/B1 U$$3825/B2 VGND VGND VPWR VPWR U$$3794/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_78_2 dadda_fa_4_78_2/A dadda_fa_4_78_2/B dadda_fa_4_78_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_79_0/CIN dadda_fa_5_78_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_115_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_48_0 dadda_fa_7_48_0/A dadda_fa_7_48_0/B dadda_fa_7_48_0/CIN VGND VGND
+ VPWR VPWR _345_/D _216_/D sky130_fd_sc_hd__fa_1
XFILLER_125_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_51_0 U$$109/X U$$242/X U$$375/X VGND VGND VPWR VPWR dadda_fa_2_52_0/B
+ dadda_fa_2_51_3/B sky130_fd_sc_hd__fa_1
XFILLER_56_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_950 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$904 U$$82/A1 U$$904/A2 U$$82/B1 U$$904/B2 VGND VGND VPWR VPWR U$$905/A sky130_fd_sc_hd__a22o_1
XU$$915 U$$915/A U$$958/A VGND VGND VPWR VPWR U$$915/X sky130_fd_sc_hd__xor2_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$926 U$$926/A1 U$$942/A2 U$$928/A1 U$$942/B2 VGND VGND VPWR VPWR U$$927/A sky130_fd_sc_hd__a22o_1
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$937 U$$937/A U$$959/A VGND VGND VPWR VPWR U$$937/X sky130_fd_sc_hd__xor2_1
XFILLER_44_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$948 U$$948/A1 U$$956/A2 U$$950/A1 U$$956/B2 VGND VGND VPWR VPWR U$$949/A sky130_fd_sc_hd__a22o_1
XU$$959 U$$959/A VGND VGND VPWR VPWR U$$959/Y sky130_fd_sc_hd__inv_1
XFILLER_16_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1109 U$$1109/A U$$1171/B VGND VGND VPWR VPWR U$$1109/X sky130_fd_sc_hd__xor2_1
XFILLER_44_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_80_2 dadda_fa_3_80_2/A dadda_fa_3_80_2/B dadda_fa_3_80_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_1/A dadda_fa_4_80_2/B sky130_fd_sc_hd__fa_1
XFILLER_113_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_998 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_73_1 dadda_fa_3_73_1/A dadda_fa_3_73_1/B dadda_fa_3_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_0/CIN dadda_fa_4_73_2/A sky130_fd_sc_hd__fa_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_50_0 dadda_fa_6_50_0/A dadda_fa_6_50_0/B dadda_fa_6_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_51_0/B dadda_fa_7_50_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_66_0 dadda_fa_3_66_0/A dadda_fa_3_66_0/B dadda_fa_3_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_0/B dadda_fa_4_66_1/CIN sky130_fd_sc_hd__fa_1
Xfanout1210 U$$989/B1 VGND VGND VPWR VPWR U$$991/A1 sky130_fd_sc_hd__buf_4
Xfanout1221 input67/X VGND VGND VPWR VPWR U$$987/B1 sky130_fd_sc_hd__buf_4
Xfanout1232 U$$4412/A1 VGND VGND VPWR VPWR U$$3314/B1 sky130_fd_sc_hd__buf_2
Xfanout1243 U$$651/B VGND VGND VPWR VPWR U$$631/B sky130_fd_sc_hd__buf_6
Xfanout1254 U$$548/A VGND VGND VPWR VPWR U$$536/B sky130_fd_sc_hd__buf_4
Xfanout1265 U$$4374/B VGND VGND VPWR VPWR U$$4368/B sky130_fd_sc_hd__buf_6
XFILLER_120_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1276 U$$4191/B VGND VGND VPWR VPWR U$$4215/B sky130_fd_sc_hd__buf_6
XFILLER_19_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1287 U$$339/B VGND VGND VPWR VPWR U$$347/B sky130_fd_sc_hd__buf_2
XU$$3001 U$$3684/B1 U$$3005/A2 U$$3551/A1 U$$3005/B2 VGND VGND VPWR VPWR U$$3002/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1298 fanout1299/X VGND VGND VPWR VPWR U$$4058/B sky130_fd_sc_hd__buf_8
XU$$3012 U$$3012/A U$$3013/A VGND VGND VPWR VPWR U$$3012/X sky130_fd_sc_hd__xor2_1
XU$$3023 U$$3023/A U$$3061/B VGND VGND VPWR VPWR U$$3023/X sky130_fd_sc_hd__xor2_1
XU$$3034 U$$979/A1 U$$3124/A2 U$$979/B1 U$$3124/B2 VGND VGND VPWR VPWR U$$3035/A sky130_fd_sc_hd__a22o_1
XU$$2300 U$$2574/A1 U$$2310/A2 U$$2576/A1 U$$2310/B2 VGND VGND VPWR VPWR U$$2301/A
+ sky130_fd_sc_hd__a22o_1
XU$$3045 U$$3045/A U$$3123/B VGND VGND VPWR VPWR U$$3045/X sky130_fd_sc_hd__xor2_1
XU$$3056 U$$3056/A1 U$$3066/A2 U$$3056/B1 U$$3066/B2 VGND VGND VPWR VPWR U$$3057/A
+ sky130_fd_sc_hd__a22o_1
XU$$2311 U$$2311/A U$$2329/A VGND VGND VPWR VPWR U$$2311/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_102_1 dadda_fa_4_102_1/A dadda_fa_4_102_1/B dadda_fa_4_102_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_103_0/B dadda_fa_5_102_1/B sky130_fd_sc_hd__fa_1
XU$$3067 U$$3067/A U$$3073/B VGND VGND VPWR VPWR U$$3067/X sky130_fd_sc_hd__xor2_1
XU$$2322 U$$3966/A1 U$$2326/A2 U$$3966/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2323/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2333 U$$2331/Y input28/X U$$2329/A U$$2332/X U$$2329/Y VGND VGND VPWR VPWR U$$2333/X
+ sky130_fd_sc_hd__a32o_2
XU$$3078 U$$612/A1 U$$3124/A2 U$$3080/A1 U$$3124/B2 VGND VGND VPWR VPWR U$$3079/A
+ sky130_fd_sc_hd__a22o_1
XU$$3089 U$$3089/A U$$3151/A VGND VGND VPWR VPWR U$$3089/X sky130_fd_sc_hd__xor2_1
XU$$2344 U$$2344/A U$$2412/B VGND VGND VPWR VPWR U$$2344/X sky130_fd_sc_hd__xor2_1
XU$$2355 U$$2629/A1 U$$2395/A2 U$$850/A1 U$$2395/B2 VGND VGND VPWR VPWR U$$2356/A
+ sky130_fd_sc_hd__a22o_1
XU$$1610 U$$1610/A U$$1626/B VGND VGND VPWR VPWR U$$1610/X sky130_fd_sc_hd__xor2_1
XU$$2366 U$$2366/A U$$2402/B VGND VGND VPWR VPWR U$$2366/X sky130_fd_sc_hd__xor2_1
XU$$1621 U$$4361/A1 U$$1621/A2 U$$4363/A1 U$$1621/B2 VGND VGND VPWR VPWR U$$1622/A
+ sky130_fd_sc_hd__a22o_1
XU$$1632 U$$1632/A U$$1644/A VGND VGND VPWR VPWR U$$1632/X sky130_fd_sc_hd__xor2_1
XFILLER_62_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2377 U$$4432/A1 U$$2413/A2 U$$872/A1 U$$2413/B2 VGND VGND VPWR VPWR U$$2378/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1643 U$$1644/A VGND VGND VPWR VPWR U$$1643/Y sky130_fd_sc_hd__inv_1
XU$$2388 U$$2388/A U$$2402/B VGND VGND VPWR VPWR U$$2388/X sky130_fd_sc_hd__xor2_1
XU$$1654 U$$3022/B1 U$$1696/A2 U$$2887/B1 U$$1696/B2 VGND VGND VPWR VPWR U$$1655/A
+ sky130_fd_sc_hd__a22o_1
XU$$2399 U$$3630/B1 U$$2445/A2 U$$3495/B1 U$$2445/B2 VGND VGND VPWR VPWR U$$2400/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1665 U$$1665/A U$$1699/B VGND VGND VPWR VPWR U$$1665/X sky130_fd_sc_hd__xor2_1
XU$$1676 U$$443/A1 U$$1702/A2 U$$3048/A1 U$$1702/B2 VGND VGND VPWR VPWR U$$1677/A
+ sky130_fd_sc_hd__a22o_1
XU$$1687 U$$1687/A U$$1697/B VGND VGND VPWR VPWR U$$1687/X sky130_fd_sc_hd__xor2_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_123_0 dadda_fa_7_123_0/A dadda_fa_7_123_0/B dadda_fa_7_123_0/CIN VGND
+ VGND VPWR VPWR _420_/D _291_/D sky130_fd_sc_hd__fa_1
XU$$1698 U$$54/A1 U$$1698/A2 U$$56/A1 U$$1698/B2 VGND VGND VPWR VPWR U$$1699/A sky130_fd_sc_hd__a22o_1
XFILLER_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_88_1 dadda_fa_5_88_1/A dadda_fa_5_88_1/B dadda_fa_5_88_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_89_0/B dadda_fa_7_88_0/A sky130_fd_sc_hd__fa_1
XFILLER_116_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$306 final_adder.U$$308/B final_adder.U$$306/B VGND VGND VPWR VPWR
+ final_adder.U$$432/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$317 final_adder.U$$316/B final_adder.U$$191/X final_adder.U$$189/X
+ VGND VGND VPWR VPWR final_adder.U$$317/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$328 final_adder.U$$330/B final_adder.U$$328/B VGND VGND VPWR VPWR
+ final_adder.U$$454/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$339 final_adder.U$$338/B final_adder.U$$213/X final_adder.U$$211/X
+ VGND VGND VPWR VPWR final_adder.U$$339/X sky130_fd_sc_hd__a21o_1
XFILLER_38_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$682_1911 VGND VGND VPWR VPWR U$$682_1911/HI U$$682/B1 sky130_fd_sc_hd__conb_1
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4280 U$$4280/A U$$4322/B VGND VGND VPWR VPWR U$$4280/X sky130_fd_sc_hd__xor2_1
XU$$4291 U$$4291/A1 U$$4295/A2 U$$4291/B1 U$$4295/B2 VGND VGND VPWR VPWR U$$4292/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3590 U$$3999/B1 U$$3604/A2 U$$4001/B1 U$$3604/B2 VGND VGND VPWR VPWR U$$3591/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_90_1 dadda_fa_4_90_1/A dadda_fa_4_90_1/B dadda_fa_4_90_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_91_0/B dadda_fa_5_90_1/B sky130_fd_sc_hd__fa_1
XFILLER_5_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_83_0 dadda_fa_4_83_0/A dadda_fa_4_83_0/B dadda_fa_4_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_84_0/A dadda_fa_5_83_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_104_3 dadda_fa_3_104_3/A dadda_fa_3_104_3/B dadda_fa_3_104_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_105_1/B dadda_fa_4_104_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_84_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_3_116_0_1945 VGND VGND VPWR VPWR dadda_ha_3_116_0/A dadda_ha_3_116_0_1945/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$851 final_adder.U$$754/X final_adder.U$$819/X final_adder.U$$755/X
+ VGND VGND VPWR VPWR final_adder.U$$851/X sky130_fd_sc_hd__a21o_1
XFILLER_29_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$701 U$$973/B1 U$$771/A2 U$$840/A1 U$$771/B2 VGND VGND VPWR VPWR U$$702/A sky130_fd_sc_hd__a22o_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$873 final_adder.U$$776/X final_adder.U$$729/X final_adder.U$$777/X
+ VGND VGND VPWR VPWR final_adder.U$$873/X sky130_fd_sc_hd__a21o_1
XU$$712 U$$712/A U$$744/B VGND VGND VPWR VPWR U$$712/X sky130_fd_sc_hd__xor2_1
XU$$723 U$$997/A1 U$$763/A2 U$$997/B1 U$$763/B2 VGND VGND VPWR VPWR U$$724/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$895 final_adder.U$$798/X final_adder.U$$381/X final_adder.U$$799/X
+ VGND VGND VPWR VPWR final_adder.U$$895/X sky130_fd_sc_hd__a21o_1
XU$$734 U$$734/A U$$768/B VGND VGND VPWR VPWR U$$734/X sky130_fd_sc_hd__xor2_1
XU$$745 U$$745/A1 U$$819/A2 U$$745/B1 U$$819/B2 VGND VGND VPWR VPWR U$$746/A sky130_fd_sc_hd__a22o_1
XU$$756 U$$756/A U$$764/B VGND VGND VPWR VPWR U$$756/X sky130_fd_sc_hd__xor2_1
XU$$767 U$$902/B1 U$$769/A2 U$$84/A1 U$$769/B2 VGND VGND VPWR VPWR U$$768/A sky130_fd_sc_hd__a22o_1
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$778 U$$778/A U$$778/B VGND VGND VPWR VPWR U$$778/X sky130_fd_sc_hd__xor2_1
XU$$789 U$$926/A1 U$$809/A2 U$$928/A1 U$$809/B2 VGND VGND VPWR VPWR U$$790/A sky130_fd_sc_hd__a22o_1
XFILLER_31_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_98_0 dadda_fa_6_98_0/A dadda_fa_6_98_0/B dadda_fa_6_98_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_99_0/B dadda_fa_7_98_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_125_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4417_1856 VGND VGND VPWR VPWR U$$4417_1856/HI U$$4417/B sky130_fd_sc_hd__conb_1
XFILLER_6_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1040 U$$4452/A1 VGND VGND VPWR VPWR U$$479/A1 sky130_fd_sc_hd__buf_4
Xfanout1051 U$$3846/B1 VGND VGND VPWR VPWR U$$971/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout1062 U$$2665/B1 VGND VGND VPWR VPWR U$$64/A1 sky130_fd_sc_hd__buf_4
XFILLER_94_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1073 U$$745/B1 VGND VGND VPWR VPWR U$$882/B1 sky130_fd_sc_hd__buf_4
Xfanout1084 U$$4444/A1 VGND VGND VPWR VPWR U$$4442/B1 sky130_fd_sc_hd__buf_4
Xfanout1095 U$$3205/B1 VGND VGND VPWR VPWR U$$56/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_40_4 dadda_fa_2_40_4/A dadda_fa_2_40_4/B dadda_fa_2_40_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_41_1/CIN dadda_fa_3_40_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_33_3 U$$1270/X U$$1403/X U$$1536/X VGND VGND VPWR VPWR dadda_fa_3_34_1/B
+ dadda_fa_3_33_3/B sky130_fd_sc_hd__fa_1
XU$$2130 U$$2130/A U$$2130/B VGND VGND VPWR VPWR U$$2130/X sky130_fd_sc_hd__xor2_1
XFILLER_63_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2141 U$$86/A1 U$$2189/A2 U$$88/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2142/A sky130_fd_sc_hd__a22o_1
XFILLER_35_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2152 U$$2152/A U$$2191/A VGND VGND VPWR VPWR U$$2152/X sky130_fd_sc_hd__xor2_1
XU$$2163 U$$2574/A1 U$$2177/A2 U$$2576/A1 U$$2177/B2 VGND VGND VPWR VPWR U$$2164/A
+ sky130_fd_sc_hd__a22o_1
XU$$2174 U$$2174/A U$$2192/A VGND VGND VPWR VPWR U$$2174/X sky130_fd_sc_hd__xor2_1
XU$$2185 U$$3966/A1 U$$2189/A2 U$$3966/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2186/A
+ sky130_fd_sc_hd__a22o_1
XU$$1440 U$$481/A1 U$$1452/A2 U$$72/A1 U$$1452/B2 VGND VGND VPWR VPWR U$$1441/A sky130_fd_sc_hd__a22o_1
XU$$1451 U$$1451/A U$$1455/B VGND VGND VPWR VPWR U$$1451/X sky130_fd_sc_hd__xor2_1
XU$$2196 U$$2194/Y input26/X U$$2192/A U$$2195/X U$$2192/Y VGND VGND VPWR VPWR U$$2196/X
+ sky130_fd_sc_hd__a32o_4
XU$$1462 U$$92/A1 U$$1504/A2 U$$94/A1 U$$1504/B2 VGND VGND VPWR VPWR U$$1463/A sky130_fd_sc_hd__a22o_1
XU$$1473 U$$1473/A U$$1475/B VGND VGND VPWR VPWR U$$1473/X sky130_fd_sc_hd__xor2_1
XU$$1484 U$$386/B1 U$$1502/A2 U$$253/A1 U$$1502/B2 VGND VGND VPWR VPWR U$$1485/A sky130_fd_sc_hd__a22o_1
XU$$1495 U$$1495/A U$$1497/B VGND VGND VPWR VPWR U$$1495/X sky130_fd_sc_hd__xor2_1
XFILLER_148_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_78_5 U$$3222/X U$$3355/X U$$3488/X VGND VGND VPWR VPWR dadda_fa_2_79_2/A
+ dadda_fa_2_78_5/A sky130_fd_sc_hd__fa_1
XFILLER_131_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$103 _399_/Q _271_/Q VGND VGND VPWR VPWR final_adder.U$$153/B1 final_adder.U$$152/B
+ sky130_fd_sc_hd__ha_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$114 _410_/Q _282_/Q VGND VGND VPWR VPWR final_adder.U$$911/B1 final_adder.U$$140/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$125 _421_/Q _293_/Q VGND VGND VPWR VPWR final_adder.U$$131/B1 final_adder.U$$130/B
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$136 final_adder.U$$136/A final_adder.U$$136/B VGND VGND VPWR VPWR
+ final_adder.U$$264/B sky130_fd_sc_hd__and2_1
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$147 final_adder.U$$146/B final_adder.U$$917/B1 final_adder.U$$147/B1
+ VGND VGND VPWR VPWR final_adder.U$$147/X sky130_fd_sc_hd__a21o_1
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$158 final_adder.U$$158/A final_adder.U$$158/B VGND VGND VPWR VPWR
+ final_adder.U$$286/B sky130_fd_sc_hd__and2_1
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$169 final_adder.U$$168/B final_adder.U$$939/B1 final_adder.U$$169/B1
+ VGND VGND VPWR VPWR final_adder.U$$169/X sky130_fd_sc_hd__a21o_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_102_0 U$$4068/X U$$4201/X U$$4334/X VGND VGND VPWR VPWR dadda_fa_4_103_0/B
+ dadda_fa_4_102_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput110 b[50] VGND VGND VPWR VPWR input110/X sky130_fd_sc_hd__clkbuf_1
Xinput121 b[60] VGND VGND VPWR VPWR input121/X sky130_fd_sc_hd__clkbuf_4
Xinput132 c[102] VGND VGND VPWR VPWR input132/X sky130_fd_sc_hd__clkbuf_4
Xinput143 c[112] VGND VGND VPWR VPWR input143/X sky130_fd_sc_hd__buf_2
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_50_3 dadda_fa_3_50_3/A dadda_fa_3_50_3/B dadda_fa_3_50_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_1/B dadda_fa_4_50_2/CIN sky130_fd_sc_hd__fa_1
Xinput154 c[122] VGND VGND VPWR VPWR input154/X sky130_fd_sc_hd__buf_2
Xdadda_fa_0_66_3 U$$1336/X U$$1469/X U$$1602/X VGND VGND VPWR VPWR dadda_fa_1_67_6/B
+ dadda_fa_1_66_8/B sky130_fd_sc_hd__fa_1
Xinput165 c[17] VGND VGND VPWR VPWR input165/X sky130_fd_sc_hd__buf_2
Xdadda_fa_3_43_2 dadda_fa_3_43_2/A dadda_fa_3_43_2/B dadda_fa_3_43_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_1/A dadda_fa_4_43_2/B sky130_fd_sc_hd__fa_1
Xinput176 c[27] VGND VGND VPWR VPWR input176/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput187 c[37] VGND VGND VPWR VPWR input187/X sky130_fd_sc_hd__buf_2
XFILLER_64_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput198 c[47] VGND VGND VPWR VPWR input198/X sky130_fd_sc_hd__dlymetal6s2s_1
Xdadda_fa_0_59_2 U$$923/X U$$1056/X U$$1189/X VGND VGND VPWR VPWR dadda_fa_1_60_7/A
+ dadda_fa_1_59_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_63_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$670 final_adder.U$$686/B final_adder.U$$670/B VGND VGND VPWR VPWR
+ final_adder.U$$782/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$681 final_adder.U$$680/B final_adder.U$$577/X final_adder.U$$561/X
+ VGND VGND VPWR VPWR final_adder.U$$681/X sky130_fd_sc_hd__a21o_1
XFILLER_45_931 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$520 U$$520/A U$$522/B VGND VGND VPWR VPWR U$$520/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_36_1 dadda_fa_3_36_1/A dadda_fa_3_36_1/B dadda_fa_3_36_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_0/CIN dadda_fa_4_36_2/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$692 final_adder.U$$708/B final_adder.U$$692/B VGND VGND VPWR VPWR
+ final_adder.U$$772/A sky130_fd_sc_hd__and2_1
XU$$531 U$$805/A1 U$$539/A2 U$$805/B1 U$$539/B2 VGND VGND VPWR VPWR U$$532/A sky130_fd_sc_hd__a22o_1
XFILLER_45_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$542 U$$542/A U$$548/A VGND VGND VPWR VPWR U$$542/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_13_0 dadda_fa_6_13_0/A dadda_fa_6_13_0/B dadda_fa_6_13_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_14_0/B dadda_fa_7_13_0/CIN sky130_fd_sc_hd__fa_1
XU$$553 U$$551/B U$$548/A U$$549/A U$$548/Y VGND VGND VPWR VPWR U$$553/X sky130_fd_sc_hd__a22o_2
Xdadda_fa_3_29_0 U$$1528/X U$$1661/X U$$1794/X VGND VGND VPWR VPWR dadda_fa_4_30_0/B
+ dadda_fa_4_29_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_17_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$564 U$$975/A1 U$$610/A2 U$$566/A1 U$$610/B2 VGND VGND VPWR VPWR U$$565/A sky130_fd_sc_hd__a22o_1
XU$$575 U$$575/A U$$639/B VGND VGND VPWR VPWR U$$575/X sky130_fd_sc_hd__xor2_1
XFILLER_60_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$586 U$$721/B1 U$$636/A2 U$$999/A1 U$$636/B2 VGND VGND VPWR VPWR U$$587/A sky130_fd_sc_hd__a22o_1
XU$$597 U$$597/A U$$631/B VGND VGND VPWR VPWR U$$597/X sky130_fd_sc_hd__xor2_1
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_95_5 input251/X dadda_fa_2_95_5/B dadda_fa_2_95_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_96_2/A dadda_fa_4_95_0/A sky130_fd_sc_hd__fa_2
XFILLER_114_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_88_4 dadda_fa_2_88_4/A dadda_fa_2_88_4/B dadda_fa_2_88_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_89_1/CIN dadda_fa_3_88_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_2_25_1 U$$456/X U$$589/X VGND VGND VPWR VPWR dadda_fa_3_26_3/A dadda_fa_4_25_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_82_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_31_0 U$$69/X U$$202/X U$$335/X VGND VGND VPWR VPWR dadda_fa_3_32_0/CIN
+ dadda_fa_3_31_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_63_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1270 U$$1270/A U$$1282/B VGND VGND VPWR VPWR U$$1270/X sky130_fd_sc_hd__xor2_1
XFILLER_51_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1281 U$$48/A1 U$$1311/A2 U$$50/A1 U$$1311/B2 VGND VGND VPWR VPWR U$$1282/A sky130_fd_sc_hd__a22o_1
XU$$1292 U$$1292/A U$$1294/B VGND VGND VPWR VPWR U$$1292/X sky130_fd_sc_hd__xor2_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_118_0 dadda_fa_5_118_0/A dadda_fa_5_118_0/B dadda_fa_5_118_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_119_0/A dadda_fa_6_118_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_164_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_83_3 U$$2567/X U$$2700/X U$$2833/X VGND VGND VPWR VPWR dadda_fa_2_84_2/CIN
+ dadda_fa_2_83_5/A sky130_fd_sc_hd__fa_1
XFILLER_117_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout800 U$$2812/B2 VGND VGND VPWR VPWR U$$2856/B2 sky130_fd_sc_hd__buf_6
Xfanout811 U$$2608/X VGND VGND VPWR VPWR U$$2679/B2 sky130_fd_sc_hd__buf_4
XFILLER_104_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_60_2 dadda_fa_4_60_2/A dadda_fa_4_60_2/B dadda_fa_4_60_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_61_0/CIN dadda_fa_5_60_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout822 U$$2445/B2 VGND VGND VPWR VPWR U$$2407/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_76_2 U$$2287/X U$$2420/X U$$2553/X VGND VGND VPWR VPWR dadda_fa_2_77_1/A
+ dadda_fa_2_76_4/A sky130_fd_sc_hd__fa_1
XFILLER_131_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout833 U$$2197/X VGND VGND VPWR VPWR U$$2282/B2 sky130_fd_sc_hd__buf_4
Xfanout844 U$$2006/B2 VGND VGND VPWR VPWR U$$1964/B2 sky130_fd_sc_hd__buf_4
Xfanout855 U$$1891/B2 VGND VGND VPWR VPWR U$$1859/B2 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_4_53_1 dadda_fa_4_53_1/A dadda_fa_4_53_1/B dadda_fa_4_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_54_0/B dadda_fa_5_53_1/B sky130_fd_sc_hd__fa_1
Xfanout866 U$$1760/B2 VGND VGND VPWR VPWR U$$1720/B2 sky130_fd_sc_hd__buf_4
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_69_1 U$$2805/X U$$2938/X U$$3071/X VGND VGND VPWR VPWR dadda_fa_2_70_0/CIN
+ dadda_fa_2_69_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_7_30_0 dadda_fa_7_30_0/A dadda_fa_7_30_0/B dadda_fa_7_30_0/CIN VGND VGND
+ VPWR VPWR _327_/D _198_/D sky130_fd_sc_hd__fa_2
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout877 U$$1625/B2 VGND VGND VPWR VPWR U$$1635/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout888 U$$1460/B2 VGND VGND VPWR VPWR U$$1426/B2 sky130_fd_sc_hd__buf_4
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_46_0 dadda_fa_4_46_0/A dadda_fa_4_46_0/B dadda_fa_4_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_47_0/A dadda_fa_5_46_1/A sky130_fd_sc_hd__fa_1
Xfanout899 U$$1238/X VGND VGND VPWR VPWR U$$1361/B2 sky130_fd_sc_hd__clkbuf_4
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_361_ _361_/CLK _361_/D VGND VGND VPWR VPWR _361_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_292_ _420_/CLK _292_/D VGND VGND VPWR VPWR _292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_98_3 dadda_fa_3_98_3/A dadda_fa_3_98_3/B dadda_fa_3_98_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_99_1/B dadda_fa_4_98_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_ha_0_72_3 U$$1747/X U$$1880/X VGND VGND VPWR VPWR dadda_fa_1_73_8/A dadda_fa_2_72_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_170_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_71_1 U$$947/X U$$1080/X U$$1213/X VGND VGND VPWR VPWR dadda_fa_1_72_7/A
+ dadda_fa_1_71_8/B sky130_fd_sc_hd__fa_1
XFILLER_110_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_64_0 U$$135/X U$$268/X U$$401/X VGND VGND VPWR VPWR dadda_fa_1_65_5/B
+ dadda_fa_1_64_7/B sky130_fd_sc_hd__fa_1
XFILLER_3_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$350 U$$487/A1 U$$352/A2 U$$487/B1 U$$352/B2 VGND VGND VPWR VPWR U$$351/A sky130_fd_sc_hd__a22o_1
XFILLER_18_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$361 U$$361/A U$$363/B VGND VGND VPWR VPWR U$$361/X sky130_fd_sc_hd__xor2_1
XFILLER_91_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$372 U$$920/A1 U$$408/A2 U$$922/A1 U$$408/B2 VGND VGND VPWR VPWR U$$373/A sky130_fd_sc_hd__a22o_1
XU$$383 U$$383/A U$$387/B VGND VGND VPWR VPWR U$$383/X sky130_fd_sc_hd__xor2_1
XU$$394 U$$805/A1 U$$406/A2 U$$805/B1 U$$406/B2 VGND VGND VPWR VPWR U$$395/A sky130_fd_sc_hd__a22o_1
XFILLER_33_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4501_1898 VGND VGND VPWR VPWR U$$4501_1898/HI U$$4501/B sky130_fd_sc_hd__conb_1
XFILLER_121_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_93_2 U$$3651/X U$$3784/X U$$3917/X VGND VGND VPWR VPWR dadda_fa_3_94_1/A
+ dadda_fa_3_93_3/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_70_1 dadda_fa_5_70_1/A dadda_fa_5_70_1/B dadda_fa_5_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_71_0/B dadda_fa_7_70_0/A sky130_fd_sc_hd__fa_1
XFILLER_99_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_86_1 U$$4169/X U$$4302/X U$$4435/X VGND VGND VPWR VPWR dadda_fa_3_87_0/CIN
+ dadda_fa_3_86_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_63_0 dadda_fa_5_63_0/A dadda_fa_5_63_0/B dadda_fa_5_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_64_0/A dadda_fa_6_63_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_79_0 dadda_fa_2_79_0/A dadda_fa_2_79_0/B dadda_fa_2_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_0/B dadda_fa_3_79_2/B sky130_fd_sc_hd__fa_1
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_62_8 dadda_fa_1_62_8/A dadda_fa_1_62_8/B dadda_fa_1_62_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_63_3/A dadda_fa_3_62_0/A sky130_fd_sc_hd__fa_2
XFILLER_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1026 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_55_7 U$$3575/X U$$3708/X input207/X VGND VGND VPWR VPWR dadda_fa_2_56_2/CIN
+ dadda_fa_2_55_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4469_1882 VGND VGND VPWR VPWR U$$4469_1882/HI U$$4469/B sky130_fd_sc_hd__conb_1
Xdadda_fa_1_48_6 U$$2497/X U$$2630/X U$$2763/X VGND VGND VPWR VPWR dadda_fa_2_49_3/A
+ dadda_fa_2_48_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_82_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_956 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_78_0 dadda_fa_7_78_0/A dadda_fa_7_78_0/B dadda_fa_7_78_0/CIN VGND VGND
+ VPWR VPWR _375_/D _246_/D sky130_fd_sc_hd__fa_1
XFILLER_151_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_81_0 U$$1232/Y U$$1366/X U$$1499/X VGND VGND VPWR VPWR dadda_fa_2_82_1/A
+ dadda_fa_2_81_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_144_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1606 U$$4508/A1 VGND VGND VPWR VPWR U$$3684/B1 sky130_fd_sc_hd__buf_4
XFILLER_160_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1617 U$$2860/B1 VGND VGND VPWR VPWR U$$4506/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout630 U$$1460/A2 VGND VGND VPWR VPWR U$$1432/A2 sky130_fd_sc_hd__buf_2
XFILLER_144_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1628 U$$940/A1 VGND VGND VPWR VPWR U$$803/A1 sky130_fd_sc_hd__buf_4
XFILLER_120_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1639 input114/X VGND VGND VPWR VPWR U$$938/A1 sky130_fd_sc_hd__buf_4
Xfanout641 U$$1311/A2 VGND VGND VPWR VPWR U$$1309/A2 sky130_fd_sc_hd__buf_4
Xfanout652 U$$1100/X VGND VGND VPWR VPWR U$$1202/A2 sky130_fd_sc_hd__buf_4
XU$$4109 U$$4110/A VGND VGND VPWR VPWR U$$4109/Y sky130_fd_sc_hd__inv_1
Xfanout663 U$$904/B2 VGND VGND VPWR VPWR U$$876/B2 sky130_fd_sc_hd__buf_4
Xfanout674 U$$819/B2 VGND VGND VPWR VPWR U$$817/B2 sky130_fd_sc_hd__buf_6
Xfanout685 U$$4309/B2 VGND VGND VPWR VPWR U$$4289/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout696 U$$416/X VGND VGND VPWR VPWR U$$543/B2 sky130_fd_sc_hd__buf_4
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3408 U$$4093/A1 U$$3418/A2 U$$4093/B1 U$$3418/B2 VGND VGND VPWR VPWR U$$3409/A
+ sky130_fd_sc_hd__a22o_1
XU$$3419 U$$3419/A U$$3424/A VGND VGND VPWR VPWR U$$3419/X sky130_fd_sc_hd__xor2_1
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2707 U$$2707/A1 U$$2707/A2 U$$2707/B1 U$$2707/B2 VGND VGND VPWR VPWR U$$2708/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2718 U$$2718/A U$$2739/A VGND VGND VPWR VPWR U$$2718/X sky130_fd_sc_hd__xor2_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2729 U$$2729/A1 U$$2737/A2 U$$950/A1 U$$2737/B2 VGND VGND VPWR VPWR U$$2730/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_413_ _421_/CLK _413_/D VGND VGND VPWR VPWR _413_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_344_ _344_/CLK _344_/D VGND VGND VPWR VPWR _344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_275_ _405_/CLK _275_/D VGND VGND VPWR VPWR _275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_80_0 dadda_fa_6_80_0/A dadda_fa_6_80_0/B dadda_fa_6_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_81_0/B dadda_fa_7_80_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_96_0 dadda_fa_3_96_0/A dadda_fa_3_96_0/B dadda_fa_3_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_0/B dadda_fa_4_96_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_127_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_58_5 dadda_fa_2_58_5/A dadda_fa_2_58_5/B dadda_fa_2_58_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_2/A dadda_fa_4_58_0/A sky130_fd_sc_hd__fa_2
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3920 U$$3920/A1 U$$3924/A2 U$$908/A1 U$$3924/B2 VGND VGND VPWR VPWR U$$3921/A
+ sky130_fd_sc_hd__a22o_1
XU$$3931 U$$3931/A U$$3949/B VGND VGND VPWR VPWR U$$3931/X sky130_fd_sc_hd__xor2_1
XFILLER_64_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3942 U$$4490/A1 U$$3948/A2 U$$4081/A1 U$$3948/B2 VGND VGND VPWR VPWR U$$3943/A
+ sky130_fd_sc_hd__a22o_1
XU$$3953 U$$3953/A U$$3965/B VGND VGND VPWR VPWR U$$3953/X sky130_fd_sc_hd__xor2_1
XU$$3964 U$$3964/A1 U$$3966/A2 U$$3966/A1 U$$3966/B2 VGND VGND VPWR VPWR U$$3965/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3975 U$$4040/B VGND VGND VPWR VPWR U$$3975/Y sky130_fd_sc_hd__inv_1
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3986 U$$3986/A U$$4026/B VGND VGND VPWR VPWR U$$3986/X sky130_fd_sc_hd__xor2_1
XU$$3997 U$$4132/B1 U$$4025/A2 U$$3999/A1 U$$4025/B2 VGND VGND VPWR VPWR U$$3998/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$180 U$$180/A U$$180/B VGND VGND VPWR VPWR U$$180/X sky130_fd_sc_hd__xor2_1
XU$$191 U$$465/A1 U$$229/A2 U$$465/B1 U$$229/B2 VGND VGND VPWR VPWR U$$192/A sky130_fd_sc_hd__a22o_1
XFILLER_33_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4499_1897 VGND VGND VPWR VPWR U$$4499_1897/HI U$$4499/B sky130_fd_sc_hd__conb_1
XFILLER_119_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput266 output266/A VGND VGND VPWR VPWR o[108] sky130_fd_sc_hd__buf_2
Xoutput277 output277/A VGND VGND VPWR VPWR o[118] sky130_fd_sc_hd__buf_2
XFILLER_142_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput288 output288/A VGND VGND VPWR VPWR o[12] sky130_fd_sc_hd__buf_2
Xoutput299 output299/A VGND VGND VPWR VPWR o[22] sky130_fd_sc_hd__buf_2
XFILLER_102_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_60_5 U$$3984/X U$$4117/X U$$4133/B VGND VGND VPWR VPWR dadda_fa_2_61_2/A
+ dadda_fa_2_60_5/A sky130_fd_sc_hd__fa_1
XFILLER_56_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_4 U$$1975/X U$$2108/X U$$2241/X VGND VGND VPWR VPWR dadda_fa_2_54_1/CIN
+ dadda_fa_2_53_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_46_3 U$$1296/X U$$1429/X U$$1562/X VGND VGND VPWR VPWR dadda_fa_2_47_2/CIN
+ dadda_fa_2_46_5/A sky130_fd_sc_hd__fa_1
XFILLER_71_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_23_2 dadda_fa_4_23_2/A dadda_fa_4_23_2/B dadda_fa_4_23_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_24_0/CIN dadda_fa_5_23_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_128_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_16_1 U$$1103/X U$$1171/B input164/X VGND VGND VPWR VPWR dadda_fa_5_17_0/B
+ dadda_fa_5_16_1/B sky130_fd_sc_hd__fa_1
XFILLER_24_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1107 final_adder.U$$172/B final_adder.U$$943/X VGND VGND VPWR VPWR
+ output366/A sky130_fd_sc_hd__xor2_1
XFILLER_165_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1118 final_adder.U$$160/A final_adder.U$$869/X VGND VGND VPWR VPWR
+ output378/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1129 final_adder.U$$150/B final_adder.U$$921/X VGND VGND VPWR VPWR
+ output263/A sky130_fd_sc_hd__xor2_1
XFILLER_20_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1403 U$$2745/A2 VGND VGND VPWR VPWR U$$2668/B sky130_fd_sc_hd__buf_6
Xfanout1414 fanout1419/X VGND VGND VPWR VPWR U$$2603/A sky130_fd_sc_hd__buf_6
XFILLER_120_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1425 U$$821/A VGND VGND VPWR VPWR U$$778/B sky130_fd_sc_hd__buf_4
XFILLER_120_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1436 fanout1438/X VGND VGND VPWR VPWR U$$2456/B sky130_fd_sc_hd__buf_6
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1447 U$$2273/B VGND VGND VPWR VPWR U$$2328/A sky130_fd_sc_hd__buf_4
Xfanout1458 U$$2007/B VGND VGND VPWR VPWR U$$1963/B sky130_fd_sc_hd__buf_6
XFILLER_47_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout460 U$$3912/A2 VGND VGND VPWR VPWR U$$3872/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout1469 U$$1882/B VGND VGND VPWR VPWR U$$1832/B sky130_fd_sc_hd__buf_4
Xfanout471 U$$3703/X VGND VGND VPWR VPWR U$$3777/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout482 U$$3658/A2 VGND VGND VPWR VPWR U$$3692/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout493 U$$3292/X VGND VGND VPWR VPWR U$$3338/A2 sky130_fd_sc_hd__buf_4
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3205 U$$602/A1 U$$3207/A2 U$$3205/B1 U$$3207/B2 VGND VGND VPWR VPWR U$$3206/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3216 U$$3216/A U$$3258/B VGND VGND VPWR VPWR U$$3216/X sky130_fd_sc_hd__xor2_1
XU$$3227 U$$3636/B1 U$$3241/A2 U$$3638/B1 U$$3241/B2 VGND VGND VPWR VPWR U$$3228/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3238 U$$3238/A U$$3242/B VGND VGND VPWR VPWR U$$3238/X sky130_fd_sc_hd__xor2_1
XFILLER_74_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3249 U$$3249/A1 U$$3251/A2 U$$3249/B1 U$$3251/B2 VGND VGND VPWR VPWR U$$3250/A
+ sky130_fd_sc_hd__a22o_1
XU$$2504 U$$447/B1 U$$2548/A2 U$$2780/A1 U$$2548/B2 VGND VGND VPWR VPWR U$$2505/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2515 U$$2515/A U$$2549/B VGND VGND VPWR VPWR U$$2515/X sky130_fd_sc_hd__xor2_1
XU$$2526 U$$3072/B1 U$$2532/A2 U$$2665/A1 U$$2532/B2 VGND VGND VPWR VPWR U$$2527/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2537 U$$2537/A U$$2603/A VGND VGND VPWR VPWR U$$2537/X sky130_fd_sc_hd__xor2_1
XFILLER_61_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1803 U$$707/A1 U$$1841/A2 U$$709/A1 U$$1841/B2 VGND VGND VPWR VPWR U$$1804/A sky130_fd_sc_hd__a22o_1
XU$$2548 U$$80/B1 U$$2548/A2 U$$3920/A1 U$$2548/B2 VGND VGND VPWR VPWR U$$2549/A sky130_fd_sc_hd__a22o_1
XU$$2559 U$$2559/A U$$2603/A VGND VGND VPWR VPWR U$$2559/X sky130_fd_sc_hd__xor2_1
XU$$1814 U$$1814/A U$$1836/B VGND VGND VPWR VPWR U$$1814/X sky130_fd_sc_hd__xor2_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1825 U$$864/B1 U$$1829/A2 U$$729/B1 U$$1829/B2 VGND VGND VPWR VPWR U$$1826/A sky130_fd_sc_hd__a22o_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1836 U$$1836/A U$$1836/B VGND VGND VPWR VPWR U$$1836/X sky130_fd_sc_hd__xor2_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1847 U$$612/B1 U$$1881/A2 U$$479/A1 U$$1881/B2 VGND VGND VPWR VPWR U$$1848/A sky130_fd_sc_hd__a22o_1
XU$$1858 U$$1858/A U$$1882/B VGND VGND VPWR VPWR U$$1858/X sky130_fd_sc_hd__xor2_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1869 U$$3376/A1 U$$1909/A2 U$$88/B1 U$$1909/B2 VGND VGND VPWR VPWR U$$1870/A sky130_fd_sc_hd__a22o_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_327_ _344_/CLK _327_/D VGND VGND VPWR VPWR _327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_258_ _258_/CLK _258_/D VGND VGND VPWR VPWR _258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_189_ _321_/CLK _189_/D VGND VGND VPWR VPWR _189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_70_4 dadda_fa_2_70_4/A dadda_fa_2_70_4/B dadda_fa_2_70_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_1/CIN dadda_fa_3_70_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_97_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_63_3 dadda_fa_2_63_3/A dadda_fa_2_63_3/B dadda_fa_2_63_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_1/B dadda_fa_3_63_3/B sky130_fd_sc_hd__fa_1
XFILLER_78_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_56_2 dadda_fa_2_56_2/A dadda_fa_2_56_2/B dadda_fa_2_56_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_1/A dadda_fa_3_56_3/A sky130_fd_sc_hd__fa_1
XU$$4440 U$$4440/A1 U$$4388/X U$$4440/B1 U$$4516/B2 VGND VGND VPWR VPWR U$$4441/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_33_1 dadda_fa_5_33_1/A dadda_fa_5_33_1/B dadda_fa_5_33_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_34_0/B dadda_fa_7_33_0/A sky130_fd_sc_hd__fa_1
XFILLER_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4451 U$$4451/A U$$4451/B VGND VGND VPWR VPWR U$$4451/X sky130_fd_sc_hd__xor2_1
XFILLER_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_49_1 dadda_fa_2_49_1/A dadda_fa_2_49_1/B dadda_fa_2_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_0/CIN dadda_fa_3_49_2/CIN sky130_fd_sc_hd__fa_1
XU$$4462 U$$4462/A1 U$$4388/X U$$4464/A1 U$$4488/B2 VGND VGND VPWR VPWR U$$4463/A
+ sky130_fd_sc_hd__a22o_1
XU$$4473 U$$4473/A U$$4473/B VGND VGND VPWR VPWR U$$4473/X sky130_fd_sc_hd__xor2_1
XU$$4484 U$$4484/A1 U$$4388/X U$$4484/B1 U$$4488/B2 VGND VGND VPWR VPWR U$$4485/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_26_0 dadda_fa_5_26_0/A dadda_fa_5_26_0/B dadda_fa_5_26_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_27_0/A dadda_fa_6_26_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_92_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3750 U$$3750/A U$$3828/B VGND VGND VPWR VPWR U$$3750/X sky130_fd_sc_hd__xor2_1
XU$$4495 U$$4495/A U$$4495/B VGND VGND VPWR VPWR U$$4495/X sky130_fd_sc_hd__xor2_1
XU$$3761 U$$4307/B1 U$$3773/A2 U$$3763/A1 U$$3773/B2 VGND VGND VPWR VPWR U$$3762/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3772 U$$3772/A U$$3774/B VGND VGND VPWR VPWR U$$3772/X sky130_fd_sc_hd__xor2_1
XFILLER_53_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3783 U$$4468/A1 U$$3829/A2 U$$4470/A1 U$$3829/B2 VGND VGND VPWR VPWR U$$3784/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3794 U$$3794/A U$$3816/B VGND VGND VPWR VPWR U$$3794/X sky130_fd_sc_hd__xor2_1
XFILLER_52_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_100_0 dadda_fa_5_100_0/A dadda_fa_5_100_0/B dadda_fa_5_100_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_101_0/A dadda_fa_6_100_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_173_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_51_1 U$$508/X U$$641/X U$$774/X VGND VGND VPWR VPWR dadda_fa_2_52_0/CIN
+ dadda_fa_2_51_3/CIN sky130_fd_sc_hd__fa_1
XU$$905 U$$905/A U$$907/B VGND VGND VPWR VPWR U$$905/X sky130_fd_sc_hd__xor2_1
XU$$916 U$$916/A1 U$$956/A2 U$$918/A1 U$$956/B2 VGND VGND VPWR VPWR U$$917/A sky130_fd_sc_hd__a22o_1
XU$$927 U$$927/A U$$959/A VGND VGND VPWR VPWR U$$927/X sky130_fd_sc_hd__xor2_1
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_44_0 U$$95/X U$$228/X U$$361/X VGND VGND VPWR VPWR dadda_fa_2_45_2/B dadda_fa_2_44_4/B
+ sky130_fd_sc_hd__fa_1
XFILLER_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$938 U$$938/A1 U$$942/A2 U$$940/A1 U$$942/B2 VGND VGND VPWR VPWR U$$939/A sky130_fd_sc_hd__a22o_1
XFILLER_44_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$949 U$$949/A U$$958/A VGND VGND VPWR VPWR U$$949/X sky130_fd_sc_hd__xor2_1
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_80_3 dadda_fa_3_80_3/A dadda_fa_3_80_3/B dadda_fa_3_80_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_1/B dadda_fa_4_80_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_125_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_73_2 dadda_fa_3_73_2/A dadda_fa_3_73_2/B dadda_fa_3_73_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_1/A dadda_fa_4_73_2/B sky130_fd_sc_hd__fa_1
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1200 U$$1088/B VGND VGND VPWR VPWR U$$1094/B sky130_fd_sc_hd__buf_6
XFILLER_79_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1211 U$$852/B1 VGND VGND VPWR VPWR U$$989/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_66_1 dadda_fa_3_66_1/A dadda_fa_3_66_1/B dadda_fa_3_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_0/CIN dadda_fa_4_66_2/A sky130_fd_sc_hd__fa_1
Xfanout1222 U$$3181/A1 VGND VGND VPWR VPWR U$$576/B1 sky130_fd_sc_hd__buf_4
Xfanout1233 input66/X VGND VGND VPWR VPWR U$$4412/A1 sky130_fd_sc_hd__buf_6
Xfanout1244 U$$651/B VGND VGND VPWR VPWR U$$637/B sky130_fd_sc_hd__buf_6
Xdadda_fa_6_43_0 dadda_fa_6_43_0/A dadda_fa_6_43_0/B dadda_fa_6_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_44_0/B dadda_fa_7_43_0/CIN sky130_fd_sc_hd__fa_1
Xfanout1255 U$$547/A VGND VGND VPWR VPWR U$$548/A sky130_fd_sc_hd__buf_4
Xdadda_fa_3_59_0 dadda_fa_3_59_0/A dadda_fa_3_59_0/B dadda_fa_3_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_0/B dadda_fa_4_59_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1266 U$$4374/B VGND VGND VPWR VPWR U$$4350/B sky130_fd_sc_hd__buf_6
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1277 U$$4191/B VGND VGND VPWR VPWR U$$4227/B sky130_fd_sc_hd__buf_4
XFILLER_19_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1288 U$$387/B VGND VGND VPWR VPWR U$$339/B sky130_fd_sc_hd__buf_4
XU$$3002 U$$3002/A U$$3004/B VGND VGND VPWR VPWR U$$3002/X sky130_fd_sc_hd__xor2_1
Xfanout1299 input55/X VGND VGND VPWR VPWR fanout1299/X sky130_fd_sc_hd__buf_4
XFILLER_115_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3013 U$$3013/A VGND VGND VPWR VPWR U$$3013/Y sky130_fd_sc_hd__inv_1
XU$$3024 U$$3296/B1 U$$3066/A2 U$$3163/A1 U$$3066/B2 VGND VGND VPWR VPWR U$$3025/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3035 U$$3035/A U$$3077/B VGND VGND VPWR VPWR U$$3035/X sky130_fd_sc_hd__xor2_1
XU$$2301 U$$2301/A U$$2301/B VGND VGND VPWR VPWR U$$2301/X sky130_fd_sc_hd__xor2_1
XFILLER_62_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3046 U$$3181/B1 U$$3124/A2 U$$3048/A1 U$$3124/B2 VGND VGND VPWR VPWR U$$3047/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3057 U$$3057/A U$$3061/B VGND VGND VPWR VPWR U$$3057/X sky130_fd_sc_hd__xor2_1
XU$$2312 U$$2312/A1 U$$2320/A2 U$$2860/B1 U$$2320/B2 VGND VGND VPWR VPWR U$$2313/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_102_2 dadda_fa_4_102_2/A dadda_fa_4_102_2/B dadda_fa_4_102_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_103_0/CIN dadda_fa_5_102_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3068 U$$4162/B1 U$$3072/A2 U$$4027/B1 U$$3072/B2 VGND VGND VPWR VPWR U$$3069/A
+ sky130_fd_sc_hd__a22o_1
XU$$2323 U$$2323/A U$$2327/B VGND VGND VPWR VPWR U$$2323/X sky130_fd_sc_hd__xor2_1
XU$$2334 U$$2332/B U$$2301/B input28/X U$$2329/Y VGND VGND VPWR VPWR U$$2334/X sky130_fd_sc_hd__a22o_2
XU$$1600 U$$1600/A U$$1608/B VGND VGND VPWR VPWR U$$1600/X sky130_fd_sc_hd__xor2_1
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3079 U$$3079/A U$$3123/B VGND VGND VPWR VPWR U$$3079/X sky130_fd_sc_hd__xor2_1
XU$$2345 U$$3850/B1 U$$2415/A2 U$$4402/A1 U$$2415/B2 VGND VGND VPWR VPWR U$$2346/A
+ sky130_fd_sc_hd__a22o_1
XU$$2356 U$$2356/A U$$2396/B VGND VGND VPWR VPWR U$$2356/X sky130_fd_sc_hd__xor2_1
XU$$1611 U$$787/B1 U$$1625/A2 U$$654/A1 U$$1625/B2 VGND VGND VPWR VPWR U$$1612/A sky130_fd_sc_hd__a22o_1
XU$$2367 U$$38/A1 U$$2415/A2 U$$40/A1 U$$2415/B2 VGND VGND VPWR VPWR U$$2368/A sky130_fd_sc_hd__a22o_1
XU$$1622 U$$1622/A U$$1626/B VGND VGND VPWR VPWR U$$1622/X sky130_fd_sc_hd__xor2_1
XU$$1633 U$$2179/B1 U$$1635/A2 U$$2183/A1 U$$1635/B2 VGND VGND VPWR VPWR U$$1634/A
+ sky130_fd_sc_hd__a22o_1
XU$$2378 U$$2378/A U$$2416/B VGND VGND VPWR VPWR U$$2378/X sky130_fd_sc_hd__xor2_1
XU$$2389 U$$3072/B1 U$$2395/A2 U$$2665/A1 U$$2395/B2 VGND VGND VPWR VPWR U$$2390/A
+ sky130_fd_sc_hd__a22o_1
XU$$1644 U$$1644/A VGND VGND VPWR VPWR U$$1644/Y sky130_fd_sc_hd__inv_1
XFILLER_62_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1655 U$$1655/A U$$1697/B VGND VGND VPWR VPWR U$$1655/X sky130_fd_sc_hd__xor2_1
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1666 U$$2897/B1 U$$1702/A2 U$$981/B1 U$$1702/B2 VGND VGND VPWR VPWR U$$1667/A
+ sky130_fd_sc_hd__a22o_1
XU$$1677 U$$1677/A U$$1703/B VGND VGND VPWR VPWR U$$1677/X sky130_fd_sc_hd__xor2_1
XU$$1688 U$$864/B1 U$$1696/A2 U$$729/B1 U$$1696/B2 VGND VGND VPWR VPWR U$$1689/A sky130_fd_sc_hd__a22o_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1699 U$$1699/A U$$1699/B VGND VGND VPWR VPWR U$$1699/X sky130_fd_sc_hd__xor2_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_116_0 dadda_fa_7_116_0/A dadda_fa_7_116_0/B dadda_fa_7_116_0/CIN VGND
+ VGND VPWR VPWR _413_/D _284_/D sky130_fd_sc_hd__fa_1
XFILLER_147_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_61_0 dadda_fa_2_61_0/A dadda_fa_2_61_0/B dadda_fa_2_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_0/B dadda_fa_3_61_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$307 final_adder.U$$306/B final_adder.U$$181/X final_adder.U$$179/X
+ VGND VGND VPWR VPWR final_adder.U$$307/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$318 final_adder.U$$320/B final_adder.U$$318/B VGND VGND VPWR VPWR
+ final_adder.U$$444/B sky130_fd_sc_hd__and2_1
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$329 final_adder.U$$328/B final_adder.U$$203/X final_adder.U$$201/X
+ VGND VGND VPWR VPWR final_adder.U$$329/X sky130_fd_sc_hd__a21o_1
XFILLER_85_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4270 U$$4270/A U$$4294/B VGND VGND VPWR VPWR U$$4270/X sky130_fd_sc_hd__xor2_1
XU$$4281 U$$4416/B1 U$$4325/A2 U$$4283/A1 U$$4325/B2 VGND VGND VPWR VPWR U$$4282/A
+ sky130_fd_sc_hd__a22o_1
XU$$4292 U$$4292/A U$$4292/B VGND VGND VPWR VPWR U$$4292/X sky130_fd_sc_hd__xor2_1
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3580 U$$3580/A1 U$$3644/A2 U$$3580/B1 U$$3644/B2 VGND VGND VPWR VPWR U$$3581/A
+ sky130_fd_sc_hd__a22o_1
XU$$3591 U$$3591/A U$$3601/B VGND VGND VPWR VPWR U$$3591/X sky130_fd_sc_hd__xor2_1
XFILLER_80_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2890 U$$2890/A U$$2926/B VGND VGND VPWR VPWR U$$2890/X sky130_fd_sc_hd__xor2_1
XFILLER_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_90_2 dadda_fa_4_90_2/A dadda_fa_4_90_2/B dadda_fa_4_90_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_91_0/CIN dadda_fa_5_90_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_174_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_83_1 dadda_fa_4_83_1/A dadda_fa_4_83_1/B dadda_fa_4_83_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_84_0/B dadda_fa_5_83_1/B sky130_fd_sc_hd__fa_1
XFILLER_135_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_60_0 dadda_fa_7_60_0/A dadda_fa_7_60_0/B dadda_fa_7_60_0/CIN VGND VGND
+ VPWR VPWR _357_/D _228_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_76_0 dadda_fa_4_76_0/A dadda_fa_4_76_0/B dadda_fa_4_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_77_0/A dadda_fa_5_76_1/A sky130_fd_sc_hd__fa_1
XFILLER_150_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$841 final_adder.U$$744/X final_adder.U$$809/X final_adder.U$$745/X
+ VGND VGND VPWR VPWR final_adder.U$$841/X sky130_fd_sc_hd__a21o_2
XFILLER_63_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$863 final_adder.U$$766/X final_adder.U$$831/X final_adder.U$$767/X
+ VGND VGND VPWR VPWR final_adder.U$$863/X sky130_fd_sc_hd__a21o_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$702 U$$702/A U$$774/B VGND VGND VPWR VPWR U$$702/X sky130_fd_sc_hd__xor2_1
XFILLER_91_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$713 U$$28/A1 U$$743/A2 U$$30/A1 U$$743/B2 VGND VGND VPWR VPWR U$$714/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$885 final_adder.U$$788/X final_adder.U$$621/X final_adder.U$$789/X
+ VGND VGND VPWR VPWR final_adder.U$$885/X sky130_fd_sc_hd__a21o_1
XU$$724 U$$724/A U$$764/B VGND VGND VPWR VPWR U$$724/X sky130_fd_sc_hd__xor2_1
XFILLER_44_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$735 U$$735/A1 U$$769/A2 U$$735/B1 U$$769/B2 VGND VGND VPWR VPWR U$$736/A sky130_fd_sc_hd__a22o_1
XU$$746 U$$746/A U$$778/B VGND VGND VPWR VPWR U$$746/X sky130_fd_sc_hd__xor2_1
XU$$757 U$$894/A1 U$$763/A2 U$$896/A1 U$$763/B2 VGND VGND VPWR VPWR U$$758/A sky130_fd_sc_hd__a22o_1
XU$$768 U$$768/A U$$768/B VGND VGND VPWR VPWR U$$768/X sky130_fd_sc_hd__xor2_1
XU$$779 U$$914/B1 U$$817/A2 U$$781/A1 U$$817/B2 VGND VGND VPWR VPWR U$$780/A sky130_fd_sc_hd__a22o_1
XFILLER_45_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$143_1788 VGND VGND VPWR VPWR U$$143_1788/HI U$$143/A1 sky130_fd_sc_hd__conb_1
XFILLER_125_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1030 U$$4315/B1 VGND VGND VPWR VPWR U$$70/A1 sky130_fd_sc_hd__buf_6
XFILLER_94_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1041 U$$4315/A1 VGND VGND VPWR VPWR U$$3628/B1 sky130_fd_sc_hd__buf_6
Xfanout1052 U$$4396/A1 VGND VGND VPWR VPWR U$$3846/B1 sky130_fd_sc_hd__buf_4
Xfanout1063 U$$2665/B1 VGND VGND VPWR VPWR U$$884/B1 sky130_fd_sc_hd__buf_2
XFILLER_94_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1074 input84/X VGND VGND VPWR VPWR U$$745/B1 sky130_fd_sc_hd__buf_6
Xfanout1085 input83/X VGND VGND VPWR VPWR U$$4444/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1096 input81/X VGND VGND VPWR VPWR U$$3205/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_40_5 dadda_fa_2_40_5/A dadda_fa_2_40_5/B dadda_fa_2_40_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_41_2/A dadda_fa_4_40_0/A sky130_fd_sc_hd__fa_2
XFILLER_94_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_33_4 U$$1669/X U$$1802/X U$$1935/X VGND VGND VPWR VPWR dadda_fa_3_34_1/CIN
+ dadda_fa_3_33_3/CIN sky130_fd_sc_hd__fa_1
XU$$2120 U$$2120/A U$$2148/B VGND VGND VPWR VPWR U$$2120/X sky130_fd_sc_hd__xor2_1
XU$$2131 U$$3636/B1 U$$2177/A2 U$$900/A1 U$$2177/B2 VGND VGND VPWR VPWR U$$2132/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2142 U$$2142/A U$$2191/A VGND VGND VPWR VPWR U$$2142/X sky130_fd_sc_hd__xor2_1
XU$$2153 U$$3249/A1 U$$2189/A2 U$$3249/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2154/A
+ sky130_fd_sc_hd__a22o_1
XU$$2164 U$$2164/A U$$2168/B VGND VGND VPWR VPWR U$$2164/X sky130_fd_sc_hd__xor2_1
XFILLER_63_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1430 U$$469/B1 U$$1460/A2 U$$884/A1 U$$1460/B2 VGND VGND VPWR VPWR U$$1431/A sky130_fd_sc_hd__a22o_1
XU$$2175 U$$2312/A1 U$$2181/A2 U$$2175/B1 U$$2181/B2 VGND VGND VPWR VPWR U$$2176/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2186 U$$2186/A U$$2186/B VGND VGND VPWR VPWR U$$2186/X sky130_fd_sc_hd__xor2_1
XU$$1441 U$$1441/A U$$1449/B VGND VGND VPWR VPWR U$$1441/X sky130_fd_sc_hd__xor2_1
XU$$2197 U$$2195/B U$$2168/B input26/X U$$2192/Y VGND VGND VPWR VPWR U$$2197/X sky130_fd_sc_hd__a22o_4
XU$$1452 U$$82/A1 U$$1452/A2 U$$82/B1 U$$1452/B2 VGND VGND VPWR VPWR U$$1453/A sky130_fd_sc_hd__a22o_1
XU$$1463 U$$1463/A U$$1475/B VGND VGND VPWR VPWR U$$1463/X sky130_fd_sc_hd__xor2_1
XFILLER_15_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1474 U$$2979/B1 U$$1504/A2 U$$928/A1 U$$1504/B2 VGND VGND VPWR VPWR U$$1475/A
+ sky130_fd_sc_hd__a22o_1
XU$$1485 U$$1485/A U$$1491/B VGND VGND VPWR VPWR U$$1485/X sky130_fd_sc_hd__xor2_1
XU$$1496 U$$2179/B1 U$$1504/A2 U$$2183/A1 U$$1504/B2 VGND VGND VPWR VPWR U$$1497/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_93_0 dadda_fa_5_93_0/A dadda_fa_5_93_0/B dadda_fa_5_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_94_0/A dadda_fa_6_93_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_78_6 U$$3621/X U$$3754/X U$$3887/X VGND VGND VPWR VPWR dadda_fa_2_79_2/B
+ dadda_fa_2_78_5/B sky130_fd_sc_hd__fa_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$104 _400_/Q _272_/Q VGND VGND VPWR VPWR final_adder.U$$921/B1 final_adder.U$$150/A
+ sky130_fd_sc_hd__ha_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$115 _411_/Q _283_/Q VGND VGND VPWR VPWR final_adder.U$$141/B1 final_adder.U$$140/B
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$126 _422_/Q _294_/Q VGND VGND VPWR VPWR final_adder.U$$899/B1 final_adder.U$$899/A1
+ sky130_fd_sc_hd__ha_2
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$137 final_adder.U$$136/B final_adder.U$$907/B1 final_adder.U$$137/B1
+ VGND VGND VPWR VPWR final_adder.U$$137/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$148 final_adder.U$$148/A final_adder.U$$148/B VGND VGND VPWR VPWR
+ final_adder.U$$276/B sky130_fd_sc_hd__and2_1
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$159 final_adder.U$$158/B final_adder.U$$929/B1 final_adder.U$$159/B1
+ VGND VGND VPWR VPWR final_adder.U$$159/X sky130_fd_sc_hd__a21o_1
XFILLER_26_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_102_1 U$$4467/X input132/X dadda_fa_3_102_1/CIN VGND VGND VPWR VPWR dadda_fa_4_103_0/CIN
+ dadda_fa_4_102_2/A sky130_fd_sc_hd__fa_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput100 b[41] VGND VGND VPWR VPWR input100/X sky130_fd_sc_hd__buf_2
XFILLER_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput111 b[51] VGND VGND VPWR VPWR input111/X sky130_fd_sc_hd__clkbuf_1
Xinput122 b[61] VGND VGND VPWR VPWR input122/X sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_6_123_0 dadda_fa_6_123_0/A dadda_fa_6_123_0/B dadda_fa_6_123_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_124_0/B dadda_fa_7_123_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput133 c[103] VGND VGND VPWR VPWR input133/X sky130_fd_sc_hd__clkbuf_4
Xinput144 c[113] VGND VGND VPWR VPWR input144/X sky130_fd_sc_hd__buf_2
Xinput155 c[123] VGND VGND VPWR VPWR input155/X sky130_fd_sc_hd__buf_2
Xdadda_fa_0_66_4 U$$1735/X U$$1868/X U$$2001/X VGND VGND VPWR VPWR dadda_fa_1_67_6/CIN
+ dadda_fa_1_66_8/CIN sky130_fd_sc_hd__fa_1
Xinput166 c[18] VGND VGND VPWR VPWR input166/X sky130_fd_sc_hd__clkbuf_4
XFILLER_102_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput177 c[28] VGND VGND VPWR VPWR input177/X sky130_fd_sc_hd__dlymetal6s2s_1
Xdadda_fa_3_43_3 dadda_fa_3_43_3/A dadda_fa_3_43_3/B dadda_fa_3_43_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_1/B dadda_fa_4_43_2/CIN sky130_fd_sc_hd__fa_1
Xinput188 c[38] VGND VGND VPWR VPWR input188/X sky130_fd_sc_hd__buf_2
XFILLER_5_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput199 c[48] VGND VGND VPWR VPWR input199/X sky130_fd_sc_hd__clkbuf_1
Xfinal_adder.U$$660 final_adder.U$$676/B final_adder.U$$660/B VGND VGND VPWR VPWR
+ final_adder.U$$772/B sky130_fd_sc_hd__and2_1
XFILLER_45_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$671 final_adder.U$$670/B final_adder.U$$567/X final_adder.U$$551/X
+ VGND VGND VPWR VPWR final_adder.U$$671/X sky130_fd_sc_hd__a21o_1
XU$$510 U$$510/A U$$522/B VGND VGND VPWR VPWR U$$510/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$682 final_adder.U$$698/B final_adder.U$$682/B VGND VGND VPWR VPWR
+ final_adder.U$$794/B sky130_fd_sc_hd__and2_1
XFILLER_29_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$521 U$$521/A1 U$$545/A2 U$$521/B1 U$$545/B2 VGND VGND VPWR VPWR U$$522/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_36_2 dadda_fa_3_36_2/A dadda_fa_3_36_2/B dadda_fa_3_36_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_1/A dadda_fa_4_36_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$693 final_adder.U$$692/B final_adder.U$$589/X final_adder.U$$573/X
+ VGND VGND VPWR VPWR final_adder.U$$693/X sky130_fd_sc_hd__a21o_1
XU$$532 U$$532/A U$$536/B VGND VGND VPWR VPWR U$$532/X sky130_fd_sc_hd__xor2_1
XFILLER_45_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$543 U$$678/B1 U$$543/A2 U$$545/A1 U$$543/B2 VGND VGND VPWR VPWR U$$544/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_29_1 U$$1927/X input178/X dadda_fa_3_29_1/CIN VGND VGND VPWR VPWR dadda_fa_4_30_0/CIN
+ dadda_fa_4_29_2/A sky130_fd_sc_hd__fa_1
XU$$554 U$$554/A1 U$$610/A2 U$$965/B1 U$$610/B2 VGND VGND VPWR VPWR U$$555/A sky130_fd_sc_hd__a22o_1
XU$$565 U$$565/A U$$607/B VGND VGND VPWR VPWR U$$565/X sky130_fd_sc_hd__xor2_1
XU$$576 U$$576/A1 U$$610/A2 U$$576/B1 U$$610/B2 VGND VGND VPWR VPWR U$$577/A sky130_fd_sc_hd__a22o_1
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$587 U$$587/A U$$637/B VGND VGND VPWR VPWR U$$587/X sky130_fd_sc_hd__xor2_1
XU$$598 U$$735/A1 U$$636/A2 U$$598/B1 U$$636/B2 VGND VGND VPWR VPWR U$$599/A sky130_fd_sc_hd__a22o_1
XFILLER_44_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_88_5 dadda_fa_2_88_5/A dadda_fa_2_88_5/B dadda_fa_2_88_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_89_2/A dadda_fa_4_88_0/A sky130_fd_sc_hd__fa_1
XFILLER_125_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_31_1 U$$468/X U$$601/X U$$734/X VGND VGND VPWR VPWR dadda_fa_3_32_1/A
+ dadda_fa_3_31_3/A sky130_fd_sc_hd__fa_1
XFILLER_74_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_24_0 U$$55/X U$$188/X U$$321/X VGND VGND VPWR VPWR dadda_fa_3_25_3/A dadda_fa_3_24_3/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_161_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1260 U$$1260/A U$$1294/B VGND VGND VPWR VPWR U$$1260/X sky130_fd_sc_hd__xor2_1
XU$$1271 U$$447/B1 U$$1309/A2 U$$314/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1272/A sky130_fd_sc_hd__a22o_1
XU$$1282 U$$1282/A U$$1282/B VGND VGND VPWR VPWR U$$1282/X sky130_fd_sc_hd__xor2_1
XFILLER_149_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1293 U$$60/A1 U$$1295/A2 U$$62/A1 U$$1295/B2 VGND VGND VPWR VPWR U$$1294/A sky130_fd_sc_hd__a22o_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_84_6 U$$3766/X U$$3899/X VGND VGND VPWR VPWR dadda_fa_2_85_4/A dadda_fa_3_84_0/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_5_118_1 dadda_fa_5_118_1/A dadda_fa_5_118_1/B dadda_ha_4_118_2/SUM VGND
+ VGND VPWR VPWR dadda_fa_6_119_0/B dadda_fa_7_118_0/A sky130_fd_sc_hd__fa_1
XFILLER_132_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_83_4 U$$2966/X U$$3099/X U$$3232/X VGND VGND VPWR VPWR dadda_fa_2_84_3/A
+ dadda_fa_2_83_5/B sky130_fd_sc_hd__fa_1
XFILLER_117_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout801 U$$2874/B2 VGND VGND VPWR VPWR U$$2872/B2 sky130_fd_sc_hd__buf_4
Xfanout812 U$$2540/B2 VGND VGND VPWR VPWR U$$2532/B2 sky130_fd_sc_hd__buf_4
XFILLER_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout823 U$$2445/B2 VGND VGND VPWR VPWR U$$2443/B2 sky130_fd_sc_hd__buf_6
XFILLER_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout834 U$$2320/B2 VGND VGND VPWR VPWR U$$2310/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_76_3 U$$2686/X U$$2819/X U$$2952/X VGND VGND VPWR VPWR dadda_fa_2_77_1/B
+ dadda_fa_2_76_4/B sky130_fd_sc_hd__fa_1
XFILLER_58_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout845 U$$2022/B2 VGND VGND VPWR VPWR U$$2006/B2 sky130_fd_sc_hd__buf_4
Xfanout856 U$$1881/B2 VGND VGND VPWR VPWR U$$1841/B2 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_4_53_2 dadda_fa_4_53_2/A dadda_fa_4_53_2/B dadda_fa_4_53_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_54_0/CIN dadda_fa_5_53_1/CIN sky130_fd_sc_hd__fa_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout867 U$$1758/B2 VGND VGND VPWR VPWR U$$1774/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_69_2 U$$3204/X U$$3337/X U$$3470/X VGND VGND VPWR VPWR dadda_fa_2_70_1/A
+ dadda_fa_2_69_4/A sky130_fd_sc_hd__fa_1
XFILLER_131_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout878 U$$1621/B2 VGND VGND VPWR VPWR U$$1625/B2 sky130_fd_sc_hd__buf_6
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_46_1 dadda_fa_4_46_1/A dadda_fa_4_46_1/B dadda_fa_4_46_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_47_0/B dadda_fa_5_46_1/B sky130_fd_sc_hd__fa_1
Xfanout889 U$$1460/B2 VGND VGND VPWR VPWR U$$1432/B2 sky130_fd_sc_hd__buf_2
XFILLER_86_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_23_0 dadda_fa_7_23_0/A dadda_fa_7_23_0/B dadda_fa_7_23_0/CIN VGND VGND
+ VPWR VPWR _320_/D _191_/D sky130_fd_sc_hd__fa_2
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_39_0 dadda_fa_4_39_0/A dadda_fa_4_39_0/B dadda_fa_4_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_40_0/A dadda_fa_5_39_1/A sky130_fd_sc_hd__fa_1
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_360_ _360_/CLK _360_/D VGND VGND VPWR VPWR _360_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_291_ _421_/CLK _291_/D VGND VGND VPWR VPWR _291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_71_2 U$$1346/X U$$1479/X U$$1612/X VGND VGND VPWR VPWR dadda_fa_1_72_7/B
+ dadda_fa_1_71_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_64_1 U$$534/X U$$667/X U$$800/X VGND VGND VPWR VPWR dadda_fa_1_65_5/CIN
+ dadda_fa_1_64_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_41_0 dadda_fa_3_41_0/A dadda_fa_3_41_0/B dadda_fa_3_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_0/B dadda_fa_4_41_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_57_0 U$$121/X U$$254/X U$$387/X VGND VGND VPWR VPWR dadda_fa_1_58_7/A
+ dadda_fa_1_57_8/B sky130_fd_sc_hd__fa_1
XFILLER_92_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$490 final_adder.U$$494/B final_adder.U$$490/B VGND VGND VPWR VPWR
+ final_adder.U$$614/B sky130_fd_sc_hd__and2_1
XU$$340 U$$749/B1 U$$340/A2 U$$616/A1 U$$340/B2 VGND VGND VPWR VPWR U$$341/A sky130_fd_sc_hd__a22o_1
XU$$351 U$$351/A U$$353/B VGND VGND VPWR VPWR U$$351/X sky130_fd_sc_hd__xor2_1
XU$$362 U$$499/A1 U$$362/A2 U$$90/A1 U$$362/B2 VGND VGND VPWR VPWR U$$363/A sky130_fd_sc_hd__a22o_1
XU$$373 U$$373/A U$$387/B VGND VGND VPWR VPWR U$$373/X sky130_fd_sc_hd__xor2_1
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$384 U$$384/A1 U$$386/A2 U$$384/B1 U$$386/B2 VGND VGND VPWR VPWR U$$385/A sky130_fd_sc_hd__a22o_1
XU$$395 U$$395/A U$$407/B VGND VGND VPWR VPWR U$$395/X sky130_fd_sc_hd__xor2_1
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_93_3 U$$4050/X U$$4183/X U$$4316/X VGND VGND VPWR VPWR dadda_fa_3_94_1/B
+ dadda_fa_3_93_3/B sky130_fd_sc_hd__fa_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_86_2 input241/X dadda_fa_2_86_2/B dadda_fa_2_86_2/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_87_1/A dadda_fa_3_86_3/A sky130_fd_sc_hd__fa_1
XFILLER_99_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_63_1 dadda_fa_5_63_1/A dadda_fa_5_63_1/B dadda_fa_5_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_64_0/B dadda_fa_7_63_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_79_1 dadda_fa_2_79_1/A dadda_fa_2_79_1/B dadda_fa_2_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_0/CIN dadda_fa_3_79_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_56_0 dadda_fa_5_56_0/A dadda_fa_5_56_0/B dadda_fa_5_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_57_0/A dadda_fa_6_56_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_55_8 dadda_fa_1_55_8/A dadda_fa_1_55_8/B dadda_fa_1_55_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_56_3/A dadda_fa_3_55_0/A sky130_fd_sc_hd__fa_1
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_102_0 dadda_fa_2_102_0/A U$$2738/X U$$2871/X VGND VGND VPWR VPWR dadda_fa_3_103_2/A
+ dadda_fa_3_102_3/A sky130_fd_sc_hd__fa_1
XFILLER_24_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1090 U$$1090/A U$$1094/B VGND VGND VPWR VPWR U$$1090/X sky130_fd_sc_hd__xor2_1
XFILLER_164_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_81_1 U$$1632/X U$$1765/X U$$1898/X VGND VGND VPWR VPWR dadda_fa_2_82_1/B
+ dadda_fa_2_81_4/A sky130_fd_sc_hd__fa_1
Xfanout1607 U$$4508/A1 VGND VGND VPWR VPWR U$$3960/A1 sky130_fd_sc_hd__buf_2
Xfanout1618 input117/X VGND VGND VPWR VPWR U$$2860/B1 sky130_fd_sc_hd__buf_6
XFILLER_160_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout620 U$$1511/X VGND VGND VPWR VPWR U$$1621/A2 sky130_fd_sc_hd__buf_8
Xdadda_fa_1_74_0 U$$1751/X U$$1884/X U$$2017/X VGND VGND VPWR VPWR dadda_fa_2_75_0/B
+ dadda_fa_2_74_3/B sky130_fd_sc_hd__fa_1
Xfanout631 U$$1480/A2 VGND VGND VPWR VPWR U$$1460/A2 sky130_fd_sc_hd__buf_4
Xfanout1629 U$$940/A1 VGND VGND VPWR VPWR U$$2310/A1 sky130_fd_sc_hd__buf_4
Xfanout642 U$$1353/A2 VGND VGND VPWR VPWR U$$1311/A2 sky130_fd_sc_hd__buf_4
XFILLER_120_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout653 U$$999/B2 VGND VGND VPWR VPWR U$$997/B2 sky130_fd_sc_hd__buf_4
XFILLER_59_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout664 U$$904/B2 VGND VGND VPWR VPWR U$$910/B2 sky130_fd_sc_hd__buf_2
Xfanout675 U$$690/X VGND VGND VPWR VPWR U$$819/B2 sky130_fd_sc_hd__buf_4
XFILLER_19_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout686 U$$4309/B2 VGND VGND VPWR VPWR U$$4381/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_74_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout697 U$$545/B2 VGND VGND VPWR VPWR U$$447/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3409 U$$3409/A U$$3411/B VGND VGND VPWR VPWR U$$3409/X sky130_fd_sc_hd__xor2_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2708 U$$2708/A U$$2708/B VGND VGND VPWR VPWR U$$2708/X sky130_fd_sc_hd__xor2_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2719 U$$4363/A1 U$$2733/A2 U$$4365/A1 U$$2733/B2 VGND VGND VPWR VPWR U$$2720/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_412_ _421_/CLK _412_/D VGND VGND VPWR VPWR _412_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_343_ _343_/CLK _343_/D VGND VGND VPWR VPWR _343_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_274_ _402_/CLK _274_/D VGND VGND VPWR VPWR _274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_96_1 dadda_fa_3_96_1/A dadda_fa_3_96_1/B dadda_fa_3_96_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_0/CIN dadda_fa_4_96_2/A sky130_fd_sc_hd__fa_1
XFILLER_170_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_73_0 dadda_fa_6_73_0/A dadda_fa_6_73_0/B dadda_fa_6_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_74_0/B dadda_fa_7_73_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_89_0 dadda_fa_3_89_0/A dadda_fa_3_89_0/B dadda_fa_3_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_0/B dadda_fa_4_89_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3910 U$$4458/A1 U$$3912/A2 U$$4049/A1 U$$3912/B2 VGND VGND VPWR VPWR U$$3911/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_118_0 dadda_fa_4_118_0/A U$$3834/X U$$3967/X VGND VGND VPWR VPWR dadda_fa_5_119_0/B
+ dadda_fa_5_118_1/A sky130_fd_sc_hd__fa_1
XU$$3921 U$$3921/A U$$3925/B VGND VGND VPWR VPWR U$$3921/X sky130_fd_sc_hd__xor2_1
XFILLER_94_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3932 U$$4478/B1 U$$3948/A2 U$$4345/A1 U$$3948/B2 VGND VGND VPWR VPWR U$$3933/A
+ sky130_fd_sc_hd__a22o_1
XU$$3943 U$$3943/A U$$3949/B VGND VGND VPWR VPWR U$$3943/X sky130_fd_sc_hd__xor2_1
XFILLER_64_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3954 U$$4365/A1 U$$3970/A2 U$$4365/B1 U$$3970/B2 VGND VGND VPWR VPWR U$$3955/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3965 U$$3965/A U$$3965/B VGND VGND VPWR VPWR U$$3965/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_5_5_0 U$$17/X U$$150/X VGND VGND VPWR VPWR dadda_fa_6_6_0/B dadda_fa_7_5_0/A
+ sky130_fd_sc_hd__ha_1
XU$$3976 U$$4110/A U$$3976/B VGND VGND VPWR VPWR U$$3976/X sky130_fd_sc_hd__and2_1
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3987 U$$4259/B1 U$$4025/A2 U$$4400/A1 U$$4025/B2 VGND VGND VPWR VPWR U$$3988/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3998 U$$3998/A U$$4026/B VGND VGND VPWR VPWR U$$3998/X sky130_fd_sc_hd__xor2_1
XU$$170 U$$170/A U$$210/B VGND VGND VPWR VPWR U$$170/X sky130_fd_sc_hd__xor2_1
XU$$181 U$$44/A1 U$$213/A2 U$$46/A1 U$$213/B2 VGND VGND VPWR VPWR U$$182/A sky130_fd_sc_hd__a22o_1
XU$$192 U$$192/A U$$230/B VGND VGND VPWR VPWR U$$192/X sky130_fd_sc_hd__xor2_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_91_0 U$$3115/X U$$3248/X U$$3381/X VGND VGND VPWR VPWR dadda_fa_3_92_0/B
+ dadda_fa_3_91_2/B sky130_fd_sc_hd__fa_1
Xoutput267 output267/A VGND VGND VPWR VPWR o[109] sky130_fd_sc_hd__buf_2
Xoutput278 output278/A VGND VGND VPWR VPWR o[119] sky130_fd_sc_hd__buf_2
Xoutput289 output289/A VGND VGND VPWR VPWR o[13] sky130_fd_sc_hd__buf_2
XFILLER_142_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_47_6 U$$2495/X U$$2628/X VGND VGND VPWR VPWR dadda_fa_2_48_3/B dadda_fa_3_47_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_101_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_60_6 input213/X dadda_fa_1_60_6/B dadda_fa_1_60_6/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_61_2/B dadda_fa_2_60_5/B sky130_fd_sc_hd__fa_2
XFILLER_68_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_53_5 U$$2374/X U$$2507/X U$$2640/X VGND VGND VPWR VPWR dadda_fa_2_54_2/A
+ dadda_fa_2_53_5/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_46_4 U$$1695/X U$$1828/X U$$1961/X VGND VGND VPWR VPWR dadda_fa_2_47_3/A
+ dadda_fa_2_46_5/B sky130_fd_sc_hd__fa_1
XFILLER_43_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_16_2 dadda_fa_4_16_2/A dadda_fa_4_16_2/B dadda_ha_3_16_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_17_0/CIN dadda_fa_5_16_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_51_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_90_0 dadda_fa_7_90_0/A dadda_fa_7_90_0/B dadda_fa_7_90_0/CIN VGND VGND
+ VPWR VPWR _387_/D _258_/D sky130_fd_sc_hd__fa_2
XFILLER_149_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1108 final_adder.U$$170/A final_adder.U$$879/X VGND VGND VPWR VPWR
+ output367/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1119 final_adder.U$$160/B final_adder.U$$931/X VGND VGND VPWR VPWR
+ output379/A sky130_fd_sc_hd__xor2_1
XFILLER_20_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1404 U$$2708/B VGND VGND VPWR VPWR U$$2740/A sky130_fd_sc_hd__buf_6
Xfanout1415 fanout1419/X VGND VGND VPWR VPWR U$$2545/B sky130_fd_sc_hd__buf_6
Xfanout1426 U$$821/A VGND VGND VPWR VPWR U$$774/B sky130_fd_sc_hd__buf_6
Xfanout1437 fanout1438/X VGND VGND VPWR VPWR U$$2465/A sky130_fd_sc_hd__buf_2
XFILLER_120_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout450 U$$4043/A2 VGND VGND VPWR VPWR U$$4025/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout1448 input27/X VGND VGND VPWR VPWR U$$2273/B sky130_fd_sc_hd__buf_6
Xfanout1459 U$$2054/A VGND VGND VPWR VPWR U$$2007/B sky130_fd_sc_hd__buf_6
Xfanout461 U$$3912/A2 VGND VGND VPWR VPWR U$$3906/A2 sky130_fd_sc_hd__buf_4
Xfanout472 U$$3703/X VGND VGND VPWR VPWR U$$3791/A2 sky130_fd_sc_hd__buf_6
XFILLER_150_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout483 U$$3566/X VGND VGND VPWR VPWR U$$3658/A2 sky130_fd_sc_hd__buf_4
Xfanout494 U$$3292/X VGND VGND VPWR VPWR U$$3340/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3206 U$$3206/A U$$3208/B VGND VGND VPWR VPWR U$$3206/X sky130_fd_sc_hd__xor2_1
XFILLER_171_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3217 U$$4450/A1 U$$3283/A2 U$$4315/A1 U$$3283/B2 VGND VGND VPWR VPWR U$$3218/A
+ sky130_fd_sc_hd__a22o_1
XU$$3228 U$$3228/A U$$3242/B VGND VGND VPWR VPWR U$$3228/X sky130_fd_sc_hd__xor2_1
XU$$3239 U$$3239/A1 U$$3241/A2 U$$3239/B1 U$$3241/B2 VGND VGND VPWR VPWR U$$3240/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2505 U$$2505/A U$$2545/B VGND VGND VPWR VPWR U$$2505/X sky130_fd_sc_hd__xor2_1
XU$$2516 U$$872/A1 U$$2546/A2 U$$874/A1 U$$2546/B2 VGND VGND VPWR VPWR U$$2517/A sky130_fd_sc_hd__a22o_1
XU$$2527 U$$2527/A U$$2529/B VGND VGND VPWR VPWR U$$2527/X sky130_fd_sc_hd__xor2_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2538 U$$3495/B1 U$$2578/A2 U$$3499/A1 U$$2578/B2 VGND VGND VPWR VPWR U$$2539/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1804 U$$1804/A U$$1836/B VGND VGND VPWR VPWR U$$1804/X sky130_fd_sc_hd__xor2_1
XFILLER_61_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2549 U$$2549/A U$$2549/B VGND VGND VPWR VPWR U$$2549/X sky130_fd_sc_hd__xor2_1
XU$$1815 U$$854/B1 U$$1831/A2 U$$3322/B1 U$$1831/B2 VGND VGND VPWR VPWR U$$1816/A
+ sky130_fd_sc_hd__a22o_1
XU$$1826 U$$1826/A U$$1828/B VGND VGND VPWR VPWR U$$1826/X sky130_fd_sc_hd__xor2_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1837 U$$741/A1 U$$1841/A2 U$$880/A1 U$$1841/B2 VGND VGND VPWR VPWR U$$1838/A sky130_fd_sc_hd__a22o_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1848 U$$1848/A U$$1854/B VGND VGND VPWR VPWR U$$1848/X sky130_fd_sc_hd__xor2_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1859 U$$900/A1 U$$1859/A2 U$$900/B1 U$$1859/B2 VGND VGND VPWR VPWR U$$1860/A sky130_fd_sc_hd__a22o_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_326_ _344_/CLK _326_/D VGND VGND VPWR VPWR _326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_257_ _386_/CLK _257_/D VGND VGND VPWR VPWR _257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_188_ _321_/CLK _188_/D VGND VGND VPWR VPWR _188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_70_5 dadda_fa_2_70_5/A dadda_fa_2_70_5/B dadda_fa_2_70_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_2/A dadda_fa_4_70_0/A sky130_fd_sc_hd__fa_1
XFILLER_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_63_4 dadda_fa_2_63_4/A dadda_fa_2_63_4/B dadda_fa_2_63_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_1/CIN dadda_fa_3_63_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_56_3 dadda_fa_2_56_3/A dadda_fa_2_56_3/B dadda_fa_2_56_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_1/B dadda_fa_3_56_3/B sky130_fd_sc_hd__fa_1
XFILLER_37_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4430 U$$4430/A1 U$$4388/X U$$4432/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4431/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4441 U$$4441/A U$$4441/B VGND VGND VPWR VPWR U$$4441/X sky130_fd_sc_hd__xor2_1
XU$$4452 U$$4452/A1 U$$4388/X U$$4454/A1 U$$4458/B2 VGND VGND VPWR VPWR U$$4453/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_49_2 dadda_fa_2_49_2/A dadda_fa_2_49_2/B dadda_fa_2_49_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_1/A dadda_fa_3_49_3/A sky130_fd_sc_hd__fa_1
XU$$4463 U$$4463/A U$$4463/B VGND VGND VPWR VPWR U$$4463/X sky130_fd_sc_hd__xor2_1
XU$$4474 U$$4474/A1 U$$4388/X U$$4474/B1 U$$4488/B2 VGND VGND VPWR VPWR U$$4475/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_26_1 dadda_fa_5_26_1/A dadda_fa_5_26_1/B dadda_fa_5_26_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_27_0/B dadda_fa_7_26_0/A sky130_fd_sc_hd__fa_2
XU$$3740 U$$3740/A U$$3740/B VGND VGND VPWR VPWR U$$3740/X sky130_fd_sc_hd__xor2_1
XU$$4485 U$$4485/A U$$4485/B VGND VGND VPWR VPWR U$$4485/X sky130_fd_sc_hd__xor2_1
XU$$3751 U$$3751/A1 U$$3829/A2 U$$3751/B1 U$$3829/B2 VGND VGND VPWR VPWR U$$3752/A
+ sky130_fd_sc_hd__a22o_1
XU$$4496 U$$4496/A1 U$$4388/X U$$4498/A1 U$$4506/B2 VGND VGND VPWR VPWR U$$4497/A
+ sky130_fd_sc_hd__a22o_1
XU$$3762 U$$3762/A U$$3774/B VGND VGND VPWR VPWR U$$3762/X sky130_fd_sc_hd__xor2_1
XFILLER_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3773 U$$3908/B1 U$$3773/A2 U$$3775/A1 U$$3773/B2 VGND VGND VPWR VPWR U$$3774/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_19_0 dadda_fa_5_19_0/A dadda_fa_5_19_0/B dadda_fa_5_19_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_20_0/A dadda_fa_6_19_0/CIN sky130_fd_sc_hd__fa_1
XU$$3784 U$$3784/A U$$3828/B VGND VGND VPWR VPWR U$$3784/X sky130_fd_sc_hd__xor2_1
XU$$3795 U$$4480/A1 U$$3825/A2 U$$4345/A1 U$$3825/B2 VGND VGND VPWR VPWR U$$3796/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_100_1 dadda_fa_5_100_1/A dadda_fa_5_100_1/B dadda_fa_5_100_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_101_0/B dadda_fa_7_100_0/A sky130_fd_sc_hd__fa_1
XFILLER_106_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_4_122_0 dadda_ha_4_122_0/A U$$4108/X VGND VGND VPWR VPWR dadda_fa_5_123_1/CIN
+ dadda_ha_4_122_0/SUM sky130_fd_sc_hd__ha_1
XFILLER_88_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_1_38_2 U$$881/X U$$1014/X VGND VGND VPWR VPWR dadda_fa_2_39_5/A dadda_fa_3_38_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_51_2 U$$907/X U$$1040/X U$$1173/X VGND VGND VPWR VPWR dadda_fa_2_52_1/A
+ dadda_fa_2_51_4/A sky130_fd_sc_hd__fa_1
XU$$906 U$$82/B1 U$$910/A2 U$$906/B1 U$$910/B2 VGND VGND VPWR VPWR U$$907/A sky130_fd_sc_hd__a22o_1
XFILLER_83_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$917 U$$917/A U$$958/A VGND VGND VPWR VPWR U$$917/X sky130_fd_sc_hd__xor2_1
XU$$928 U$$928/A1 U$$942/A2 U$$930/A1 U$$942/B2 VGND VGND VPWR VPWR U$$929/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_44_1 U$$494/X U$$627/X U$$760/X VGND VGND VPWR VPWR dadda_fa_2_45_2/CIN
+ dadda_fa_2_44_4/CIN sky130_fd_sc_hd__fa_1
XU$$939 U$$939/A U$$943/B VGND VGND VPWR VPWR U$$939/X sky130_fd_sc_hd__xor2_1
XFILLER_83_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_21_0 input170/X dadda_fa_4_21_0/B dadda_fa_4_21_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_5_22_0/A dadda_fa_5_21_1/A sky130_fd_sc_hd__fa_1
XFILLER_37_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_37_0 U$$81/X U$$214/X U$$347/X VGND VGND VPWR VPWR dadda_fa_2_38_4/CIN
+ dadda_fa_2_37_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_73_3 dadda_fa_3_73_3/A dadda_fa_3_73_3/B dadda_fa_3_73_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_1/B dadda_fa_4_73_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1201 input7/X VGND VGND VPWR VPWR U$$1088/B sky130_fd_sc_hd__buf_4
Xdadda_fa_3_66_2 dadda_fa_3_66_2/A dadda_fa_3_66_2/B dadda_fa_3_66_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_1/A dadda_fa_4_66_2/B sky130_fd_sc_hd__fa_1
Xfanout1212 U$$854/A1 VGND VGND VPWR VPWR U$$852/B1 sky130_fd_sc_hd__buf_4
XFILLER_79_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1223 U$$3181/A1 VGND VGND VPWR VPWR U$$30/A1 sky130_fd_sc_hd__buf_4
Xfanout1234 U$$3981/A1 VGND VGND VPWR VPWR U$$3022/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1245 U$$685/A VGND VGND VPWR VPWR U$$669/B sky130_fd_sc_hd__buf_4
XFILLER_78_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_59_1 dadda_fa_3_59_1/A dadda_fa_3_59_1/B dadda_fa_3_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_0/CIN dadda_fa_4_59_2/A sky130_fd_sc_hd__fa_1
Xfanout1256 U$$522/B VGND VGND VPWR VPWR U$$448/B sky130_fd_sc_hd__buf_4
Xfanout1267 U$$4374/B VGND VGND VPWR VPWR U$$4360/B sky130_fd_sc_hd__buf_4
Xfanout1278 fanout1279/X VGND VGND VPWR VPWR U$$4191/B sky130_fd_sc_hd__buf_8
Xdadda_fa_6_36_0 dadda_fa_6_36_0/A dadda_fa_6_36_0/B dadda_fa_6_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_37_0/B dadda_fa_7_36_0/CIN sky130_fd_sc_hd__fa_1
Xfanout1289 input56/X VGND VGND VPWR VPWR U$$387/B sky130_fd_sc_hd__buf_8
XU$$3003 U$$3551/A1 U$$3005/A2 U$$3416/A1 U$$3005/B2 VGND VGND VPWR VPWR U$$3004/A
+ sky130_fd_sc_hd__a22o_1
XU$$3014 U$$3014/A VGND VGND VPWR VPWR U$$3014/Y sky130_fd_sc_hd__inv_1
XU$$3025 U$$3025/A U$$3061/B VGND VGND VPWR VPWR U$$3025/X sky130_fd_sc_hd__xor2_1
XU$$3036 U$$979/B1 U$$3122/A2 U$$3447/B1 U$$3122/B2 VGND VGND VPWR VPWR U$$3037/A
+ sky130_fd_sc_hd__a22o_1
XU$$2302 U$$2576/A1 U$$2310/A2 U$$2576/B1 U$$2310/B2 VGND VGND VPWR VPWR U$$2303/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3047 U$$3047/A U$$3077/B VGND VGND VPWR VPWR U$$3047/X sky130_fd_sc_hd__xor2_1
XU$$3058 U$$4428/A1 U$$3066/A2 U$$4430/A1 U$$3066/B2 VGND VGND VPWR VPWR U$$3059/A
+ sky130_fd_sc_hd__a22o_1
XU$$2313 U$$2313/A U$$2328/A VGND VGND VPWR VPWR U$$2313/X sky130_fd_sc_hd__xor2_1
XFILLER_35_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3069 U$$3069/A U$$3073/B VGND VGND VPWR VPWR U$$3069/X sky130_fd_sc_hd__xor2_1
XU$$2324 U$$954/A1 U$$2326/A2 U$$956/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2325/A sky130_fd_sc_hd__a22o_1
XU$$2335 U$$2335/A1 U$$2415/A2 U$$967/A1 U$$2415/B2 VGND VGND VPWR VPWR U$$2336/A
+ sky130_fd_sc_hd__a22o_1
XU$$1601 U$$94/A1 U$$1641/A2 U$$96/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1602/A sky130_fd_sc_hd__a22o_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2346 U$$2346/A U$$2412/B VGND VGND VPWR VPWR U$$2346/X sky130_fd_sc_hd__xor2_1
XU$$2357 U$$2631/A1 U$$2395/A2 U$$2631/B1 U$$2395/B2 VGND VGND VPWR VPWR U$$2358/A
+ sky130_fd_sc_hd__a22o_1
XU$$1612 U$$1612/A U$$1626/B VGND VGND VPWR VPWR U$$1612/X sky130_fd_sc_hd__xor2_1
XU$$1623 U$$253/A1 U$$1625/A2 U$$253/B1 U$$1625/B2 VGND VGND VPWR VPWR U$$1624/A sky130_fd_sc_hd__a22o_1
XU$$2368 U$$2368/A U$$2412/B VGND VGND VPWR VPWR U$$2368/X sky130_fd_sc_hd__xor2_1
XU$$1634 U$$1634/A U$$1644/A VGND VGND VPWR VPWR U$$1634/X sky130_fd_sc_hd__xor2_1
XU$$2379 U$$50/A1 U$$2413/A2 U$$50/B1 U$$2413/B2 VGND VGND VPWR VPWR U$$2380/A sky130_fd_sc_hd__a22o_1
XU$$1645 input17/X VGND VGND VPWR VPWR U$$1647/B sky130_fd_sc_hd__inv_1
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1656 U$$2887/B1 U$$1696/A2 U$$2754/A1 U$$1696/B2 VGND VGND VPWR VPWR U$$1657/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1667 U$$1667/A U$$1703/B VGND VGND VPWR VPWR U$$1667/X sky130_fd_sc_hd__xor2_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1678 U$$34/A1 U$$1702/A2 U$$36/A1 U$$1702/B2 VGND VGND VPWR VPWR U$$1679/A sky130_fd_sc_hd__a22o_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1689 U$$1689/A U$$1697/B VGND VGND VPWR VPWR U$$1689/X sky130_fd_sc_hd__xor2_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_309_ _328_/CLK _309_/D VGND VGND VPWR VPWR _309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_109_0 dadda_fa_7_109_0/A dadda_fa_7_109_0/B dadda_fa_7_109_0/CIN VGND
+ VGND VPWR VPWR _406_/D _277_/D sky130_fd_sc_hd__fa_1
XFILLER_162_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_61_1 dadda_fa_2_61_1/A dadda_fa_2_61_1/B dadda_fa_2_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_0/CIN dadda_fa_3_61_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$308 final_adder.U$$310/B final_adder.U$$308/B VGND VGND VPWR VPWR
+ final_adder.U$$434/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$319 final_adder.U$$318/B final_adder.U$$193/X final_adder.U$$191/X
+ VGND VGND VPWR VPWR final_adder.U$$319/X sky130_fd_sc_hd__a21o_1
XFILLER_84_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_54_0 dadda_fa_2_54_0/A dadda_fa_2_54_0/B dadda_fa_2_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_0/B dadda_fa_3_54_2/B sky130_fd_sc_hd__fa_1
XFILLER_84_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4260 U$$4260/A U$$4292/B VGND VGND VPWR VPWR U$$4260/X sky130_fd_sc_hd__xor2_1
XFILLER_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4271 U$$4271/A1 U$$4289/A2 U$$985/A1 U$$4289/B2 VGND VGND VPWR VPWR U$$4272/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4282 U$$4282/A U$$4322/B VGND VGND VPWR VPWR U$$4282/X sky130_fd_sc_hd__xor2_1
XU$$4293 U$$4430/A1 U$$4295/A2 U$$4432/A1 U$$4295/B2 VGND VGND VPWR VPWR U$$4294/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3570 U$$3979/B1 U$$3656/A2 U$$3846/A1 U$$3656/B2 VGND VGND VPWR VPWR U$$3571/A
+ sky130_fd_sc_hd__a22o_1
XU$$3581 U$$3581/A U$$3601/B VGND VGND VPWR VPWR U$$3581/X sky130_fd_sc_hd__xor2_1
XU$$3592 U$$4001/B1 U$$3604/A2 U$$854/A1 U$$3604/B2 VGND VGND VPWR VPWR U$$3593/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2880 U$$3014/A U$$2880/B VGND VGND VPWR VPWR U$$2880/X sky130_fd_sc_hd__and2_1
Xdadda_fa_5_8_0 U$$289/X U$$422/X U$$555/X VGND VGND VPWR VPWR dadda_fa_6_9_0/A dadda_fa_6_8_0/CIN
+ sky130_fd_sc_hd__fa_1
XU$$2891 U$$3163/B1 U$$2929/A2 U$$2891/B1 U$$2929/B2 VGND VGND VPWR VPWR U$$2892/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_83_2 dadda_fa_4_83_2/A dadda_fa_4_83_2/B dadda_fa_4_83_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_84_0/CIN dadda_fa_5_83_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_150_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_76_1 dadda_fa_4_76_1/A dadda_fa_4_76_1/B dadda_fa_4_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_77_0/B dadda_fa_5_76_1/B sky130_fd_sc_hd__fa_1
XFILLER_150_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_53_0 dadda_fa_7_53_0/A dadda_fa_7_53_0/B dadda_fa_7_53_0/CIN VGND VGND
+ VPWR VPWR _350_/D _221_/D sky130_fd_sc_hd__fa_1
XFILLER_115_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_69_0 dadda_fa_4_69_0/A dadda_fa_4_69_0/B dadda_fa_4_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_70_0/A dadda_fa_5_69_1/A sky130_fd_sc_hd__fa_1
XFILLER_103_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$831 final_adder.U$$798/A final_adder.U$$381/X final_adder.U$$719/X
+ VGND VGND VPWR VPWR final_adder.U$$831/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$853 final_adder.U$$756/X final_adder.U$$821/X final_adder.U$$757/X
+ VGND VGND VPWR VPWR final_adder.U$$853/X sky130_fd_sc_hd__a21o_1
XFILLER_152_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$703 U$$840/A1 U$$771/A2 U$$840/B1 U$$771/B2 VGND VGND VPWR VPWR U$$704/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$875 final_adder.U$$778/X final_adder.U$$731/X final_adder.U$$779/X
+ VGND VGND VPWR VPWR final_adder.U$$875/X sky130_fd_sc_hd__a21o_1
XFILLER_28_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$714 U$$714/A U$$744/B VGND VGND VPWR VPWR U$$714/X sky130_fd_sc_hd__xor2_1
XU$$725 U$$997/B1 U$$763/A2 U$$864/A1 U$$763/B2 VGND VGND VPWR VPWR U$$726/A sky130_fd_sc_hd__a22o_1
XFILLER_84_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$897 final_adder.U$$800/X final_adder.U$$255/X final_adder.U$$801/X
+ VGND VGND VPWR VPWR final_adder.U$$897/X sky130_fd_sc_hd__a21o_1
XU$$736 U$$736/A U$$768/B VGND VGND VPWR VPWR U$$736/X sky130_fd_sc_hd__xor2_1
XU$$747 U$$882/B1 U$$771/A2 U$$747/B1 U$$771/B2 VGND VGND VPWR VPWR U$$748/A sky130_fd_sc_hd__a22o_1
XFILLER_83_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$758 U$$758/A U$$764/B VGND VGND VPWR VPWR U$$758/X sky130_fd_sc_hd__xor2_1
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$769 U$$84/A1 U$$769/A2 U$$86/A1 U$$769/B2 VGND VGND VPWR VPWR U$$770/A sky130_fd_sc_hd__a22o_1
XFILLER_45_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_71_0 dadda_fa_3_71_0/A dadda_fa_3_71_0/B dadda_fa_3_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_0/B dadda_fa_4_71_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1020 U$$1195/B VGND VGND VPWR VPWR U$$1163/B sky130_fd_sc_hd__buf_6
Xfanout1031 U$$479/B1 VGND VGND VPWR VPWR U$$481/A1 sky130_fd_sc_hd__buf_4
Xfanout1042 U$$4315/A1 VGND VGND VPWR VPWR U$$4176/B1 sky130_fd_sc_hd__buf_4
XFILLER_94_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1053 input87/X VGND VGND VPWR VPWR U$$4396/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1064 input85/X VGND VGND VPWR VPWR U$$2665/B1 sky130_fd_sc_hd__buf_4
Xfanout1075 U$$4309/A1 VGND VGND VPWR VPWR U$$4307/B1 sky130_fd_sc_hd__buf_4
Xfanout1086 U$$56/B1 VGND VGND VPWR VPWR U$$58/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1097 U$$878/A1 VGND VGND VPWR VPWR U$$741/A1 sky130_fd_sc_hd__buf_4
XFILLER_47_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2110 U$$2110/A U$$2148/B VGND VGND VPWR VPWR U$$2110/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_100_0 dadda_fa_4_100_0/A dadda_fa_4_100_0/B dadda_fa_4_100_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_101_0/A dadda_fa_5_100_1/A sky130_fd_sc_hd__fa_1
XU$$2121 U$$66/A1 U$$2139/A2 U$$68/A1 U$$2139/B2 VGND VGND VPWR VPWR U$$2122/A sky130_fd_sc_hd__a22o_1
XFILLER_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2132 U$$2132/A U$$2140/B VGND VGND VPWR VPWR U$$2132/X sky130_fd_sc_hd__xor2_1
XU$$2143 U$$3650/A1 U$$2189/A2 U$$3650/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2144/A
+ sky130_fd_sc_hd__a22o_1
XU$$2154 U$$2154/A U$$2191/A VGND VGND VPWR VPWR U$$2154/X sky130_fd_sc_hd__xor2_1
XU$$1420 U$$596/B1 U$$1426/A2 U$$598/B1 U$$1426/B2 VGND VGND VPWR VPWR U$$1421/A sky130_fd_sc_hd__a22o_1
XU$$2165 U$$2576/A1 U$$2177/A2 U$$2576/B1 U$$2177/B2 VGND VGND VPWR VPWR U$$2166/A
+ sky130_fd_sc_hd__a22o_1
XU$$1431 U$$1431/A U$$1461/B VGND VGND VPWR VPWR U$$1431/X sky130_fd_sc_hd__xor2_1
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2176 U$$2176/A U$$2192/A VGND VGND VPWR VPWR U$$2176/X sky130_fd_sc_hd__xor2_1
XU$$1442 U$$72/A1 U$$1452/A2 U$$74/A1 U$$1452/B2 VGND VGND VPWR VPWR U$$1443/A sky130_fd_sc_hd__a22o_1
XU$$2187 U$$3966/B1 U$$2189/A2 U$$3833/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2188/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2198 U$$2198/A1 U$$2254/A2 U$$2748/A1 U$$2254/B2 VGND VGND VPWR VPWR U$$2199/A
+ sky130_fd_sc_hd__a22o_1
XU$$1453 U$$1453/A U$$1455/B VGND VGND VPWR VPWR U$$1453/X sky130_fd_sc_hd__xor2_1
XU$$1464 U$$3106/B1 U$$1504/A2 U$$2973/A1 U$$1504/B2 VGND VGND VPWR VPWR U$$1465/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1475 U$$1475/A U$$1475/B VGND VGND VPWR VPWR U$$1475/X sky130_fd_sc_hd__xor2_1
XU$$1486 U$$251/B1 U$$1502/A2 U$$253/B1 U$$1502/B2 VGND VGND VPWR VPWR U$$1487/A sky130_fd_sc_hd__a22o_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1497 U$$1497/A U$$1497/B VGND VGND VPWR VPWR U$$1497/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_93_1 dadda_fa_5_93_1/A dadda_fa_5_93_1/B dadda_fa_5_93_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_94_0/B dadda_fa_7_93_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_86_0 dadda_fa_5_86_0/A dadda_fa_5_86_0/B dadda_fa_5_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_87_0/A dadda_fa_6_86_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_78_7 U$$4020/X U$$4153/X U$$4286/X VGND VGND VPWR VPWR dadda_fa_2_79_2/CIN
+ dadda_fa_2_78_5/CIN sky130_fd_sc_hd__fa_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$105 _401_/Q _273_/Q VGND VGND VPWR VPWR final_adder.U$$151/B1 final_adder.U$$150/B
+ sky130_fd_sc_hd__ha_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$116 _412_/Q _284_/Q VGND VGND VPWR VPWR final_adder.U$$909/B1 final_adder.U$$138/A
+ sky130_fd_sc_hd__ha_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$127 _423_/Q _295_/Q VGND VGND VPWR VPWR final_adder.U$$127/COUT final_adder.U$$1151/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$138 final_adder.U$$138/A final_adder.U$$138/B VGND VGND VPWR VPWR
+ final_adder.U$$266/B sky130_fd_sc_hd__and2_1
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$149 final_adder.U$$148/B final_adder.U$$919/B1 final_adder.U$$149/B1
+ VGND VGND VPWR VPWR final_adder.U$$149/X sky130_fd_sc_hd__a21o_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4090 U$$4090/A U$$4098/B VGND VGND VPWR VPWR U$$4090/X sky130_fd_sc_hd__xor2_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_102_2 dadda_fa_3_102_2/A dadda_fa_3_102_2/B dadda_fa_3_102_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_103_1/A dadda_fa_4_102_2/B sky130_fd_sc_hd__fa_1
XFILLER_147_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_927 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput101 b[42] VGND VGND VPWR VPWR input101/X sky130_fd_sc_hd__buf_2
Xinput112 b[52] VGND VGND VPWR VPWR input112/X sky130_fd_sc_hd__clkbuf_1
Xinput123 b[62] VGND VGND VPWR VPWR input123/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput134 c[104] VGND VGND VPWR VPWR input134/X sky130_fd_sc_hd__clkbuf_4
Xinput145 c[114] VGND VGND VPWR VPWR input145/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_0_66_5 U$$2134/X U$$2267/X U$$2400/X VGND VGND VPWR VPWR dadda_fa_1_67_7/A
+ dadda_fa_2_66_0/A sky130_fd_sc_hd__fa_1
Xinput156 c[124] VGND VGND VPWR VPWR input156/X sky130_fd_sc_hd__clkbuf_2
Xinput167 c[19] VGND VGND VPWR VPWR input167/X sky130_fd_sc_hd__buf_2
Xdadda_fa_6_116_0 dadda_fa_6_116_0/A dadda_fa_6_116_0/B dadda_fa_6_116_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_117_0/B dadda_fa_7_116_0/CIN sky130_fd_sc_hd__fa_1
Xinput178 c[29] VGND VGND VPWR VPWR input178/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput189 c[39] VGND VGND VPWR VPWR input189/X sky130_fd_sc_hd__buf_2
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$650 final_adder.U$$666/B final_adder.U$$650/B VGND VGND VPWR VPWR
+ final_adder.U$$762/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$661 final_adder.U$$660/B final_adder.U$$557/X final_adder.U$$541/X
+ VGND VGND VPWR VPWR final_adder.U$$661/X sky130_fd_sc_hd__a21o_1
XU$$500 U$$500/A U$$536/B VGND VGND VPWR VPWR U$$500/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$672 final_adder.U$$688/B final_adder.U$$672/B VGND VGND VPWR VPWR
+ final_adder.U$$784/B sky130_fd_sc_hd__and2_1
XFILLER_17_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$511 U$$783/B1 U$$545/A2 U$$650/A1 U$$545/B2 VGND VGND VPWR VPWR U$$512/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_36_3 dadda_fa_3_36_3/A dadda_fa_3_36_3/B dadda_fa_3_36_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_1/B dadda_fa_4_36_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$683 final_adder.U$$682/B final_adder.U$$579/X final_adder.U$$563/X
+ VGND VGND VPWR VPWR final_adder.U$$683/X sky130_fd_sc_hd__a21o_1
XU$$522 U$$522/A U$$522/B VGND VGND VPWR VPWR U$$522/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$694 final_adder.U$$710/B final_adder.U$$694/B VGND VGND VPWR VPWR
+ final_adder.U$$774/A sky130_fd_sc_hd__and2_1
XFILLER_29_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$533 U$$805/B1 U$$539/A2 U$$672/A1 U$$539/B2 VGND VGND VPWR VPWR U$$534/A sky130_fd_sc_hd__a22o_1
XFILLER_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$544 U$$544/A U$$548/A VGND VGND VPWR VPWR U$$544/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$555 U$$555/A U$$607/B VGND VGND VPWR VPWR U$$555/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_29_2 dadda_fa_3_29_2/A dadda_fa_3_29_2/B dadda_fa_3_29_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_30_1/A dadda_fa_4_29_2/B sky130_fd_sc_hd__fa_1
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$566 U$$566/A1 U$$610/A2 U$$20/A1 U$$610/B2 VGND VGND VPWR VPWR U$$567/A sky130_fd_sc_hd__a22o_1
XFILLER_45_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$577 U$$577/A U$$607/B VGND VGND VPWR VPWR U$$577/X sky130_fd_sc_hd__xor2_1
XU$$588 U$$997/B1 U$$630/A2 U$$864/A1 U$$630/B2 VGND VGND VPWR VPWR U$$589/A sky130_fd_sc_hd__a22o_1
XFILLER_112_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$599 U$$599/A U$$637/B VGND VGND VPWR VPWR U$$599/X sky130_fd_sc_hd__xor2_1
XFILLER_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_31_2 U$$867/X U$$1000/X U$$1133/X VGND VGND VPWR VPWR dadda_fa_3_32_1/B
+ dadda_fa_3_31_3/B sky130_fd_sc_hd__fa_1
XU$$1250 U$$1250/A U$$1282/B VGND VGND VPWR VPWR U$$1250/X sky130_fd_sc_hd__xor2_1
XU$$1261 U$$850/A1 U$$1295/A2 U$$989/A1 U$$1295/B2 VGND VGND VPWR VPWR U$$1262/A sky130_fd_sc_hd__a22o_1
XU$$1272 U$$1272/A U$$1278/B VGND VGND VPWR VPWR U$$1272/X sky130_fd_sc_hd__xor2_1
XFILLER_50_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1283 U$$735/A1 U$$1327/A2 U$$52/A1 U$$1327/B2 VGND VGND VPWR VPWR U$$1284/A sky130_fd_sc_hd__a22o_1
XU$$1294 U$$1294/A U$$1294/B VGND VGND VPWR VPWR U$$1294/X sky130_fd_sc_hd__xor2_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_5 U$$3365/X U$$3498/X U$$3631/X VGND VGND VPWR VPWR dadda_fa_2_84_3/B
+ dadda_fa_2_83_5/CIN sky130_fd_sc_hd__fa_1
Xfanout802 U$$2812/B2 VGND VGND VPWR VPWR U$$2874/B2 sky130_fd_sc_hd__buf_6
XFILLER_89_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout813 fanout820/X VGND VGND VPWR VPWR U$$2540/B2 sky130_fd_sc_hd__buf_6
Xfanout824 U$$2334/X VGND VGND VPWR VPWR U$$2445/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_76_4 U$$3085/X U$$3218/X U$$3351/X VGND VGND VPWR VPWR dadda_fa_2_77_1/CIN
+ dadda_fa_2_76_4/CIN sky130_fd_sc_hd__fa_1
Xfanout835 U$$2320/B2 VGND VGND VPWR VPWR U$$2326/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_98_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout846 U$$2014/B2 VGND VGND VPWR VPWR U$$1986/B2 sky130_fd_sc_hd__buf_4
Xfanout857 U$$1891/B2 VGND VGND VPWR VPWR U$$1881/B2 sky130_fd_sc_hd__clkbuf_8
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout868 U$$1758/B2 VGND VGND VPWR VPWR U$$1778/B2 sky130_fd_sc_hd__clkbuf_4
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_3 U$$3603/X U$$3736/X U$$3869/X VGND VGND VPWR VPWR dadda_fa_2_70_1/B
+ dadda_fa_2_69_4/B sky130_fd_sc_hd__fa_1
XFILLER_97_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout879 U$$1512/X VGND VGND VPWR VPWR U$$1621/B2 sky130_fd_sc_hd__buf_8
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_46_2 dadda_fa_4_46_2/A dadda_fa_4_46_2/B dadda_fa_4_46_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_47_0/CIN dadda_fa_5_46_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_39_1 dadda_fa_4_39_1/A dadda_fa_4_39_1/B dadda_fa_4_39_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_40_0/B dadda_fa_5_39_1/B sky130_fd_sc_hd__fa_1
XFILLER_100_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_16_0 dadda_fa_7_16_0/A dadda_fa_7_16_0/B dadda_fa_7_16_0/CIN VGND VGND
+ VPWR VPWR _313_/D _184_/D sky130_fd_sc_hd__fa_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_290_ _421_/CLK _290_/D VGND VGND VPWR VPWR _290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_58_3 U$$1320/X U$$1453/X VGND VGND VPWR VPWR dadda_fa_1_59_7/CIN dadda_fa_2_58_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_71_3 U$$1745/X U$$1878/X U$$2011/X VGND VGND VPWR VPWR dadda_fa_1_72_7/CIN
+ dadda_fa_2_71_0/A sky130_fd_sc_hd__fa_1
XFILLER_110_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_64_2 U$$933/X U$$1066/X U$$1199/X VGND VGND VPWR VPWR dadda_fa_1_65_6/A
+ dadda_fa_1_64_8/A sky130_fd_sc_hd__fa_1
XFILLER_67_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_41_1 dadda_fa_3_41_1/A dadda_fa_3_41_1/B dadda_fa_3_41_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_0/CIN dadda_fa_4_41_2/A sky130_fd_sc_hd__fa_1
XFILLER_18_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_57_1 U$$520/X U$$653/X U$$786/X VGND VGND VPWR VPWR dadda_fa_1_58_7/B
+ dadda_fa_1_57_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_92_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$480 final_adder.U$$484/B final_adder.U$$480/B VGND VGND VPWR VPWR
+ final_adder.U$$604/B sky130_fd_sc_hd__and2_1
Xdadda_fa_3_34_0 dadda_fa_3_34_0/A dadda_fa_3_34_0/B dadda_fa_3_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_0/B dadda_fa_4_34_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$491 final_adder.U$$490/B final_adder.U$$369/X final_adder.U$$365/X
+ VGND VGND VPWR VPWR final_adder.U$$491/X sky130_fd_sc_hd__a21o_1
XU$$330 U$$465/B1 U$$362/A2 U$$58/A1 U$$362/B2 VGND VGND VPWR VPWR U$$331/A sky130_fd_sc_hd__a22o_1
XFILLER_18_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$341 U$$341/A U$$341/B VGND VGND VPWR VPWR U$$341/X sky130_fd_sc_hd__xor2_1
XU$$352 U$$487/B1 U$$352/A2 U$$902/A1 U$$352/B2 VGND VGND VPWR VPWR U$$353/A sky130_fd_sc_hd__a22o_1
XU$$363 U$$363/A U$$363/B VGND VGND VPWR VPWR U$$363/X sky130_fd_sc_hd__xor2_1
XU$$374 U$$920/B1 U$$386/A2 U$$787/A1 U$$386/B2 VGND VGND VPWR VPWR U$$375/A sky130_fd_sc_hd__a22o_1
XU$$385 U$$385/A U$$387/B VGND VGND VPWR VPWR U$$385/X sky130_fd_sc_hd__xor2_1
XU$$396 U$$805/B1 U$$406/A2 U$$672/A1 U$$406/B2 VGND VGND VPWR VPWR U$$397/A sky130_fd_sc_hd__a22o_1
XFILLER_44_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_93_4 U$$4449/X input249/X dadda_fa_2_93_4/CIN VGND VGND VPWR VPWR dadda_fa_3_94_1/CIN
+ dadda_fa_3_93_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_86_3 dadda_fa_2_86_3/A dadda_fa_2_86_3/B dadda_fa_2_86_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_87_1/B dadda_fa_3_86_3/B sky130_fd_sc_hd__fa_1
XFILLER_99_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_79_2 dadda_fa_2_79_2/A dadda_fa_2_79_2/B dadda_fa_2_79_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_1/A dadda_fa_3_79_3/A sky130_fd_sc_hd__fa_1
XFILLER_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_56_1 dadda_fa_5_56_1/A dadda_fa_5_56_1/B dadda_fa_5_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_57_0/B dadda_fa_7_56_0/A sky130_fd_sc_hd__fa_1
XFILLER_68_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_49_0 dadda_fa_5_49_0/A dadda_fa_5_49_0/B dadda_fa_5_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_50_0/A dadda_fa_6_49_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_2_23_0 U$$53/X U$$186/X VGND VGND VPWR VPWR dadda_fa_3_24_3/B dadda_fa_4_23_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_55_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_102_1 U$$3004/X U$$3137/X U$$3270/X VGND VGND VPWR VPWR dadda_fa_3_103_2/B
+ dadda_fa_3_102_3/B sky130_fd_sc_hd__fa_1
XFILLER_50_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1080 U$$1080/A U$$1094/B VGND VGND VPWR VPWR U$$1080/X sky130_fd_sc_hd__xor2_1
XU$$1091 U$$406/A1 U$$1093/A2 U$$406/B1 U$$1093/B2 VGND VGND VPWR VPWR U$$1092/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_123_0 U$$4109/Y U$$4243/X U$$4376/X VGND VGND VPWR VPWR dadda_fa_6_124_0/A
+ dadda_fa_6_123_0/CIN sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_30_clk _388_/CLK VGND VGND VPWR VPWR _258_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_81_2 U$$2031/X U$$2164/X U$$2297/X VGND VGND VPWR VPWR dadda_fa_2_82_1/CIN
+ dadda_fa_2_81_4/B sky130_fd_sc_hd__fa_1
XFILLER_104_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1608 U$$2862/B1 VGND VGND VPWR VPWR U$$4508/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout610 U$$1760/A2 VGND VGND VPWR VPWR U$$1758/A2 sky130_fd_sc_hd__buf_6
Xfanout621 U$$259/A2 VGND VGND VPWR VPWR U$$229/A2 sky130_fd_sc_hd__buf_4
Xfanout1619 U$$942/A1 VGND VGND VPWR VPWR U$$805/A1 sky130_fd_sc_hd__buf_6
XFILLER_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_74_1 U$$2150/X U$$2283/X U$$2416/X VGND VGND VPWR VPWR dadda_fa_2_75_0/CIN
+ dadda_fa_2_74_3/CIN sky130_fd_sc_hd__fa_1
Xfanout632 U$$1452/A2 VGND VGND VPWR VPWR U$$1414/A2 sky130_fd_sc_hd__buf_4
Xfanout643 U$$1353/A2 VGND VGND VPWR VPWR U$$1359/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout654 U$$1075/B2 VGND VGND VPWR VPWR U$$999/B2 sky130_fd_sc_hd__buf_6
XFILLER_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_51_0 dadda_fa_4_51_0/A dadda_fa_4_51_0/B dadda_fa_4_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_52_0/A dadda_fa_5_51_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_67_0 U$$2535/X U$$2668/X U$$2801/X VGND VGND VPWR VPWR dadda_fa_2_68_0/B
+ dadda_fa_2_67_3/B sky130_fd_sc_hd__fa_1
Xfanout665 U$$952/B2 VGND VGND VPWR VPWR U$$904/B2 sky130_fd_sc_hd__buf_4
XFILLER_101_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout676 U$$676/B2 VGND VGND VPWR VPWR U$$630/B2 sky130_fd_sc_hd__buf_4
XFILLER_59_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout687 U$$4369/B2 VGND VGND VPWR VPWR U$$4373/B2 sky130_fd_sc_hd__buf_4
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout698 U$$505/B2 VGND VGND VPWR VPWR U$$479/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2709 U$$2844/B1 U$$2711/A2 U$$2711/A1 U$$2711/B2 VGND VGND VPWR VPWR U$$2710/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_411_ _416_/CLK _411_/D VGND VGND VPWR VPWR _411_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_969 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_342_ _342_/CLK _342_/D VGND VGND VPWR VPWR _342_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_273_ _402_/CLK _273_/D VGND VGND VPWR VPWR _273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_clk _370_/CLK VGND VGND VPWR VPWR _415_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_96_2 dadda_fa_3_96_2/A dadda_fa_3_96_2/B dadda_fa_3_96_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_1/A dadda_fa_4_96_2/B sky130_fd_sc_hd__fa_1
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_89_1 dadda_fa_3_89_1/A dadda_fa_3_89_1/B dadda_fa_3_89_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_0/CIN dadda_fa_4_89_2/A sky130_fd_sc_hd__fa_1
XFILLER_135_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_66_0 dadda_fa_6_66_0/A dadda_fa_6_66_0/B dadda_fa_6_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_67_0/B dadda_fa_7_66_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3900 U$$4174/A1 U$$3906/A2 U$$4176/A1 U$$3906/B2 VGND VGND VPWR VPWR U$$3901/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3911 U$$3911/A U$$3973/A VGND VGND VPWR VPWR U$$3911/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_118_1 U$$4100/X U$$4233/X U$$4366/X VGND VGND VPWR VPWR dadda_fa_5_119_0/CIN
+ dadda_fa_5_118_1/B sky130_fd_sc_hd__fa_1
XU$$3922 U$$4196/A1 U$$3924/A2 U$$4196/B1 U$$3924/B2 VGND VGND VPWR VPWR U$$3923/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3933 U$$3933/A U$$3949/B VGND VGND VPWR VPWR U$$3933/X sky130_fd_sc_hd__xor2_1
XU$$3944 U$$4081/A1 U$$3948/A2 U$$4081/B1 U$$3948/B2 VGND VGND VPWR VPWR U$$3945/A
+ sky130_fd_sc_hd__a22o_1
XU$$3955 U$$3955/A U$$3965/B VGND VGND VPWR VPWR U$$3955/X sky130_fd_sc_hd__xor2_1
XU$$3966 U$$3966/A1 U$$3966/A2 U$$3966/B1 U$$3966/B2 VGND VGND VPWR VPWR U$$3967/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3977 U$$3975/Y input54/X U$$3973/A U$$3976/X U$$3973/Y VGND VGND VPWR VPWR U$$3977/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3988 U$$3988/A U$$4026/B VGND VGND VPWR VPWR U$$3988/X sky130_fd_sc_hd__xor2_1
XU$$160 U$$160/A U$$182/B VGND VGND VPWR VPWR U$$160/X sky130_fd_sc_hd__xor2_1
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3999 U$$3999/A1 U$$4025/A2 U$$3999/B1 U$$4025/B2 VGND VGND VPWR VPWR U$$4000/A
+ sky130_fd_sc_hd__a22o_1
XU$$171 U$$34/A1 U$$207/A2 U$$36/A1 U$$207/B2 VGND VGND VPWR VPWR U$$172/A sky130_fd_sc_hd__a22o_1
XU$$182 U$$182/A U$$182/B VGND VGND VPWR VPWR U$$182/X sky130_fd_sc_hd__xor2_1
XU$$193 U$$465/B1 U$$229/A2 U$$58/A1 U$$229/B2 VGND VGND VPWR VPWR U$$194/A sky130_fd_sc_hd__a22o_1
XFILLER_72_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_985 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_clk _370_/CLK VGND VGND VPWR VPWR _375_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_118_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_91_1 U$$3514/X U$$3647/X U$$3780/X VGND VGND VPWR VPWR dadda_fa_3_92_0/CIN
+ dadda_fa_3_91_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_173_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_84_0 U$$4032/X U$$4165/X U$$4298/X VGND VGND VPWR VPWR dadda_fa_3_85_0/B
+ dadda_fa_3_84_2/B sky130_fd_sc_hd__fa_1
Xoutput257 output257/A VGND VGND VPWR VPWR o[0] sky130_fd_sc_hd__buf_2
Xoutput268 output268/A VGND VGND VPWR VPWR o[10] sky130_fd_sc_hd__buf_2
Xoutput279 output279/A VGND VGND VPWR VPWR o[11] sky130_fd_sc_hd__buf_2
XFILLER_59_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_60_7 dadda_fa_1_60_7/A dadda_fa_1_60_7/B dadda_fa_1_60_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_61_2/CIN dadda_fa_2_60_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_6 U$$2773/X U$$2906/X U$$3039/X VGND VGND VPWR VPWR dadda_fa_2_54_2/B
+ dadda_fa_2_53_5/B sky130_fd_sc_hd__fa_1
XFILLER_83_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_46_5 U$$2094/X U$$2227/X U$$2360/X VGND VGND VPWR VPWR dadda_fa_2_47_3/B
+ dadda_fa_2_46_5/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_7_5_0 dadda_fa_7_5_0/A dadda_fa_7_5_0/B dadda_fa_7_5_0/CIN VGND VGND VPWR
+ VPWR _302_/D _173_/D sky130_fd_sc_hd__fa_1
XFILLER_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1109 final_adder.U$$170/B final_adder.U$$941/X VGND VGND VPWR VPWR
+ output368/A sky130_fd_sc_hd__xor2_1
XFILLER_164_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_83_0 dadda_fa_7_83_0/A dadda_fa_7_83_0/B dadda_fa_7_83_0/CIN VGND VGND
+ VPWR VPWR _380_/D _251_/D sky130_fd_sc_hd__fa_2
Xdadda_fa_4_99_0 dadda_fa_4_99_0/A dadda_fa_4_99_0/B dadda_fa_4_99_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_100_0/A dadda_fa_5_99_1/A sky130_fd_sc_hd__fa_1
XFILLER_109_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1405 U$$2745/A2 VGND VGND VPWR VPWR U$$2708/B sky130_fd_sc_hd__buf_6
Xfanout1416 fanout1419/X VGND VGND VPWR VPWR U$$2549/B sky130_fd_sc_hd__buf_4
Xfanout1427 U$$821/A VGND VGND VPWR VPWR U$$820/B sky130_fd_sc_hd__buf_6
Xfanout440 U$$4114/X VGND VGND VPWR VPWR U$$4190/A2 sky130_fd_sc_hd__buf_6
Xfanout1438 input29/X VGND VGND VPWR VPWR fanout1438/X sky130_fd_sc_hd__buf_6
Xfanout1449 U$$2130/B VGND VGND VPWR VPWR U$$2096/B sky130_fd_sc_hd__buf_6
Xfanout451 U$$4043/A2 VGND VGND VPWR VPWR U$$4005/A2 sky130_fd_sc_hd__buf_2
XFILLER_120_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout462 U$$3840/X VGND VGND VPWR VPWR U$$3912/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout473 U$$3833/A2 VGND VGND VPWR VPWR U$$3829/A2 sky130_fd_sc_hd__buf_4
XFILLER_19_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout484 U$$3473/A2 VGND VGND VPWR VPWR U$$3471/A2 sky130_fd_sc_hd__buf_6
XFILLER_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout495 U$$3378/A2 VGND VGND VPWR VPWR U$$3372/A2 sky130_fd_sc_hd__buf_4
XFILLER_59_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3207 U$$878/A1 U$$3207/A2 U$$878/B1 U$$3207/B2 VGND VGND VPWR VPWR U$$3208/A sky130_fd_sc_hd__a22o_1
XU$$3218 U$$3218/A U$$3284/B VGND VGND VPWR VPWR U$$3218/X sky130_fd_sc_hd__xor2_1
XU$$3229 U$$3638/B1 U$$3241/A2 U$$3503/B1 U$$3241/B2 VGND VGND VPWR VPWR U$$3230/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2506 U$$2780/A1 U$$2548/A2 U$$2780/B1 U$$2548/B2 VGND VGND VPWR VPWR U$$2507/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2517 U$$2517/A U$$2545/B VGND VGND VPWR VPWR U$$2517/X sky130_fd_sc_hd__xor2_1
XU$$2528 U$$2665/A1 U$$2540/A2 U$$2665/B1 U$$2540/B2 VGND VGND VPWR VPWR U$$2529/A
+ sky130_fd_sc_hd__a22o_1
XU$$2539 U$$2539/A U$$2603/A VGND VGND VPWR VPWR U$$2539/X sky130_fd_sc_hd__xor2_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1805 U$$24/A1 U$$1841/A2 U$$26/A1 U$$1841/B2 VGND VGND VPWR VPWR U$$1806/A sky130_fd_sc_hd__a22o_1
XU$$1816 U$$1816/A U$$1832/B VGND VGND VPWR VPWR U$$1816/X sky130_fd_sc_hd__xor2_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1827 U$$729/B1 U$$1829/A2 U$$2925/A1 U$$1829/B2 VGND VGND VPWR VPWR U$$1828/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1838 U$$1838/A U$$1854/B VGND VGND VPWR VPWR U$$1838/X sky130_fd_sc_hd__xor2_1
XFILLER_42_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1849 U$$479/A1 U$$1881/A2 U$$479/B1 U$$1881/B2 VGND VGND VPWR VPWR U$$1850/A sky130_fd_sc_hd__a22o_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ _344_/CLK _325_/D VGND VGND VPWR VPWR _325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_972 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_256_ _258_/CLK _256_/D VGND VGND VPWR VPWR _256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_187_ _321_/CLK _187_/D VGND VGND VPWR VPWR _187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_63_5 dadda_fa_2_63_5/A dadda_fa_2_63_5/B dadda_fa_2_63_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_2/A dadda_fa_4_63_0/A sky130_fd_sc_hd__fa_2
XFILLER_97_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_1_clk _201_/CLK VGND VGND VPWR VPWR _338_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4420 input70/X U$$4388/X U$$4420/B1 U$$4428/B2 VGND VGND VPWR VPWR U$$4421/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_56_4 dadda_fa_2_56_4/A dadda_fa_2_56_4/B dadda_fa_2_56_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_1/CIN dadda_fa_3_56_3/CIN sky130_fd_sc_hd__fa_1
XU$$4431 U$$4431/A U$$4431/B VGND VGND VPWR VPWR U$$4431/X sky130_fd_sc_hd__xor2_1
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4442 U$$4442/A1 U$$4388/X U$$4442/B1 U$$4508/B2 VGND VGND VPWR VPWR U$$4443/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4453 U$$4453/A U$$4453/B VGND VGND VPWR VPWR U$$4453/X sky130_fd_sc_hd__xor2_1
XFILLER_38_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_49_3 dadda_fa_2_49_3/A dadda_fa_2_49_3/B dadda_fa_2_49_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_1/B dadda_fa_3_49_3/B sky130_fd_sc_hd__fa_1
XU$$4464 U$$4464/A1 U$$4388/X U$$4464/B1 U$$4492/B2 VGND VGND VPWR VPWR U$$4465/A
+ sky130_fd_sc_hd__a22o_1
XU$$3730 U$$3730/A U$$3734/B VGND VGND VPWR VPWR U$$3730/X sky130_fd_sc_hd__xor2_1
XFILLER_64_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4475 U$$4475/A U$$4475/B VGND VGND VPWR VPWR U$$4475/X sky130_fd_sc_hd__xor2_1
XU$$3741 U$$4152/A1 U$$3791/A2 U$$4152/B1 U$$3791/B2 VGND VGND VPWR VPWR U$$3742/A
+ sky130_fd_sc_hd__a22o_1
XU$$4486 U$$4486/A1 U$$4388/X U$$4486/B1 U$$4506/B2 VGND VGND VPWR VPWR U$$4487/A
+ sky130_fd_sc_hd__a22o_1
XU$$3752 U$$3752/A U$$3828/B VGND VGND VPWR VPWR U$$3752/X sky130_fd_sc_hd__xor2_1
XU$$4497 U$$4497/A U$$4497/B VGND VGND VPWR VPWR U$$4497/X sky130_fd_sc_hd__xor2_1
XU$$3763 U$$3763/A1 U$$3773/A2 U$$4176/A1 U$$3773/B2 VGND VGND VPWR VPWR U$$3764/A
+ sky130_fd_sc_hd__a22o_1
XU$$3774 U$$3774/A U$$3774/B VGND VGND VPWR VPWR U$$3774/X sky130_fd_sc_hd__xor2_1
XFILLER_52_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3785 U$$4196/A1 U$$3825/A2 U$$4196/B1 U$$3825/B2 VGND VGND VPWR VPWR U$$3786/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_19_1 dadda_fa_5_19_1/A dadda_fa_5_19_1/B dadda_fa_5_19_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_20_0/B dadda_fa_7_19_0/A sky130_fd_sc_hd__fa_1
XU$$3796 U$$3796/A U$$3816/B VGND VGND VPWR VPWR U$$3796/X sky130_fd_sc_hd__xor2_1
XFILLER_80_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_51_3 U$$1306/X U$$1439/X U$$1572/X VGND VGND VPWR VPWR dadda_fa_2_52_1/B
+ dadda_fa_2_51_4/B sky130_fd_sc_hd__fa_1
XFILLER_28_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$907 U$$907/A U$$907/B VGND VGND VPWR VPWR U$$907/X sky130_fd_sc_hd__xor2_1
XU$$918 U$$918/A1 U$$956/A2 U$$920/A1 U$$956/B2 VGND VGND VPWR VPWR U$$919/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_44_2 U$$893/X U$$1026/X U$$1159/X VGND VGND VPWR VPWR dadda_fa_2_45_3/A
+ dadda_fa_2_44_5/A sky130_fd_sc_hd__fa_1
XU$$929 U$$929/A U$$959/A VGND VGND VPWR VPWR U$$929/X sky130_fd_sc_hd__xor2_1
XFILLER_44_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_21_1 dadda_fa_4_21_1/A dadda_fa_4_21_1/B dadda_fa_4_21_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_22_0/B dadda_fa_5_21_1/B sky130_fd_sc_hd__fa_1
XFILLER_71_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_14_0 U$$301/X U$$434/X U$$567/X VGND VGND VPWR VPWR dadda_fa_5_15_0/A
+ dadda_fa_5_14_1/A sky130_fd_sc_hd__fa_1
XFILLER_169_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1202 U$$856/A1 VGND VGND VPWR VPWR U$$993/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_66_3 dadda_fa_3_66_3/A dadda_fa_3_66_3/B dadda_fa_3_66_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_1/B dadda_fa_4_66_2/CIN sky130_fd_sc_hd__fa_1
Xfanout1213 input68/X VGND VGND VPWR VPWR U$$854/A1 sky130_fd_sc_hd__buf_6
XFILLER_120_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1224 U$$4414/A1 VGND VGND VPWR VPWR U$$3181/A1 sky130_fd_sc_hd__buf_2
Xfanout1235 U$$3981/A1 VGND VGND VPWR VPWR U$$2748/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1246 U$$651/B VGND VGND VPWR VPWR U$$685/A sky130_fd_sc_hd__buf_4
XFILLER_66_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_59_2 dadda_fa_3_59_2/A dadda_fa_3_59_2/B dadda_fa_3_59_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_1/A dadda_fa_4_59_2/B sky130_fd_sc_hd__fa_1
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1257 U$$506/B VGND VGND VPWR VPWR U$$480/B sky130_fd_sc_hd__clkbuf_4
Xfanout1268 U$$4322/B VGND VGND VPWR VPWR U$$4374/B sky130_fd_sc_hd__clkbuf_4
Xfanout1279 input58/X VGND VGND VPWR VPWR fanout1279/X sky130_fd_sc_hd__buf_4
XFILLER_59_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3004 U$$3004/A U$$3004/B VGND VGND VPWR VPWR U$$3004/X sky130_fd_sc_hd__xor2_1
XFILLER_75_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3015 input39/X VGND VGND VPWR VPWR U$$3017/B sky130_fd_sc_hd__inv_1
XFILLER_75_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_29_0 dadda_fa_6_29_0/A dadda_fa_6_29_0/B dadda_fa_6_29_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_30_0/B dadda_fa_7_29_0/CIN sky130_fd_sc_hd__fa_1
XU$$3026 U$$3163/A1 U$$3066/A2 U$$3163/B1 U$$3066/B2 VGND VGND VPWR VPWR U$$3027/A
+ sky130_fd_sc_hd__a22o_1
XU$$3037 U$$3037/A U$$3077/B VGND VGND VPWR VPWR U$$3037/X sky130_fd_sc_hd__xor2_1
XU$$2303 U$$2303/A U$$2329/A VGND VGND VPWR VPWR U$$2303/X sky130_fd_sc_hd__xor2_1
XU$$3048 U$$3048/A1 U$$3124/A2 U$$3048/B1 U$$3124/B2 VGND VGND VPWR VPWR U$$3049/A
+ sky130_fd_sc_hd__a22o_1
XU$$3059 U$$3059/A U$$3061/B VGND VGND VPWR VPWR U$$3059/X sky130_fd_sc_hd__xor2_1
XFILLER_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2314 U$$4367/B1 U$$2320/A2 U$$4234/A1 U$$2320/B2 VGND VGND VPWR VPWR U$$2315/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2325 U$$2325/A U$$2327/B VGND VGND VPWR VPWR U$$2325/X sky130_fd_sc_hd__xor2_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2336 U$$2336/A U$$2412/B VGND VGND VPWR VPWR U$$2336/X sky130_fd_sc_hd__xor2_1
XU$$1602 U$$1602/A U$$1608/B VGND VGND VPWR VPWR U$$1602/X sky130_fd_sc_hd__xor2_1
XU$$2347 U$$4402/A1 U$$2407/A2 U$$4404/A1 U$$2407/B2 VGND VGND VPWR VPWR U$$2348/A
+ sky130_fd_sc_hd__a22o_1
XU$$2358 U$$2358/A U$$2396/B VGND VGND VPWR VPWR U$$2358/X sky130_fd_sc_hd__xor2_1
XU$$1613 U$$654/A1 U$$1625/A2 U$$654/B1 U$$1625/B2 VGND VGND VPWR VPWR U$$1614/A sky130_fd_sc_hd__a22o_1
XU$$1624 U$$1624/A U$$1626/B VGND VGND VPWR VPWR U$$1624/X sky130_fd_sc_hd__xor2_1
XU$$2369 U$$314/A1 U$$2413/A2 U$$42/A1 U$$2413/B2 VGND VGND VPWR VPWR U$$2370/A sky130_fd_sc_hd__a22o_1
XU$$1635 U$$2183/A1 U$$1635/A2 U$$4512/B1 U$$1635/B2 VGND VGND VPWR VPWR U$$1636/A
+ sky130_fd_sc_hd__a22o_1
XU$$1646 U$$1777/B VGND VGND VPWR VPWR U$$1646/Y sky130_fd_sc_hd__inv_1
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1657 U$$1657/A U$$1697/B VGND VGND VPWR VPWR U$$1657/X sky130_fd_sc_hd__xor2_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1668 U$$709/A1 U$$1702/A2 U$$709/B1 U$$1702/B2 VGND VGND VPWR VPWR U$$1669/A sky130_fd_sc_hd__a22o_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1679 U$$1679/A U$$1703/B VGND VGND VPWR VPWR U$$1679/X sky130_fd_sc_hd__xor2_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_308_ _328_/CLK _308_/D VGND VGND VPWR VPWR _308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_239_ _368_/CLK _239_/D VGND VGND VPWR VPWR _239_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4433_1864 VGND VGND VPWR VPWR U$$4433_1864/HI U$$4433/B sky130_fd_sc_hd__conb_1
Xdadda_fa_2_61_2 dadda_fa_2_61_2/A dadda_fa_2_61_2/B dadda_fa_2_61_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_1/A dadda_fa_3_61_3/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$309 final_adder.U$$308/B final_adder.U$$183/X final_adder.U$$181/X
+ VGND VGND VPWR VPWR final_adder.U$$309/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_2_54_1 dadda_fa_2_54_1/A dadda_fa_2_54_1/B dadda_fa_2_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_0/CIN dadda_fa_3_54_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_942 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_31_0 dadda_fa_5_31_0/A dadda_fa_5_31_0/B dadda_fa_5_31_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_32_0/A dadda_fa_6_31_0/CIN sky130_fd_sc_hd__fa_1
XU$$4509_1902 VGND VGND VPWR VPWR U$$4509_1902/HI U$$4509/B sky130_fd_sc_hd__conb_1
Xdadda_fa_2_47_0 U$$2761/X U$$2894/X U$$3027/X VGND VGND VPWR VPWR dadda_fa_3_48_0/B
+ dadda_fa_3_47_2/B sky130_fd_sc_hd__fa_1
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4250 U$$4383/A U$$4250/B VGND VGND VPWR VPWR U$$4250/X sky130_fd_sc_hd__and2_1
XU$$4261 U$$4398/A1 U$$4295/A2 U$$4400/A1 U$$4295/B2 VGND VGND VPWR VPWR U$$4262/A
+ sky130_fd_sc_hd__a22o_1
XU$$4272 U$$4272/A U$$4294/B VGND VGND VPWR VPWR U$$4272/X sky130_fd_sc_hd__xor2_1
XU$$4283 U$$4283/A1 U$$4373/A2 U$$4422/A1 U$$4373/B2 VGND VGND VPWR VPWR U$$4284/A
+ sky130_fd_sc_hd__a22o_1
XU$$4294 U$$4294/A U$$4294/B VGND VGND VPWR VPWR U$$4294/X sky130_fd_sc_hd__xor2_1
XFILLER_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3560 U$$3560/A U$$3561/A VGND VGND VPWR VPWR U$$3560/X sky130_fd_sc_hd__xor2_1
XFILLER_81_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3571 U$$3571/A U$$3615/B VGND VGND VPWR VPWR U$$3571/X sky130_fd_sc_hd__xor2_1
XFILLER_25_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3582 U$$4265/B1 U$$3644/A2 U$$4132/A1 U$$3644/B2 VGND VGND VPWR VPWR U$$3583/A
+ sky130_fd_sc_hd__a22o_1
XU$$3593 U$$3593/A U$$3601/B VGND VGND VPWR VPWR U$$3593/X sky130_fd_sc_hd__xor2_1
XFILLER_81_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2870 U$$3692/A1 U$$2872/A2 U$$3418/B1 U$$2872/B2 VGND VGND VPWR VPWR U$$2871/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_8_1 U$$607/B input245/X dadda_ha_4_8_0/SUM VGND VGND VPWR VPWR dadda_fa_6_9_0/B
+ dadda_fa_7_8_0/A sky130_fd_sc_hd__fa_1
XFILLER_52_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2881 U$$2879/Y input37/X U$$2877/A U$$2880/X U$$2877/Y VGND VGND VPWR VPWR U$$2881/X
+ sky130_fd_sc_hd__a32o_4
XU$$2892 U$$2892/A U$$2926/B VGND VGND VPWR VPWR U$$2892/X sky130_fd_sc_hd__xor2_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_76_2 dadda_fa_4_76_2/A dadda_fa_4_76_2/B dadda_fa_4_76_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_77_0/CIN dadda_fa_5_76_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_69_1 dadda_fa_4_69_1/A dadda_fa_4_69_1/B dadda_fa_4_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_70_0/B dadda_fa_5_69_1/B sky130_fd_sc_hd__fa_1
XFILLER_88_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_46_0 dadda_fa_7_46_0/A dadda_fa_7_46_0/B dadda_fa_7_46_0/CIN VGND VGND
+ VPWR VPWR _343_/D _214_/D sky130_fd_sc_hd__fa_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$821 final_adder.U$$788/A final_adder.U$$621/X final_adder.U$$709/X
+ VGND VGND VPWR VPWR final_adder.U$$821/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$843 final_adder.U$$746/X final_adder.U$$811/X final_adder.U$$747/X
+ VGND VGND VPWR VPWR final_adder.U$$843/X sky130_fd_sc_hd__a21o_2
XFILLER_21_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$865 final_adder.U$$768/X final_adder.U$$833/X final_adder.U$$769/X
+ VGND VGND VPWR VPWR final_adder.U$$865/X sky130_fd_sc_hd__a21o_1
XU$$704 U$$704/A U$$774/B VGND VGND VPWR VPWR U$$704/X sky130_fd_sc_hd__xor2_1
XU$$715 U$$987/B1 U$$771/A2 U$$852/B1 U$$771/B2 VGND VGND VPWR VPWR U$$716/A sky130_fd_sc_hd__a22o_1
XFILLER_56_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$887 final_adder.U$$790/X final_adder.U$$623/X final_adder.U$$791/X
+ VGND VGND VPWR VPWR final_adder.U$$887/X sky130_fd_sc_hd__a21o_1
XFILLER_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$726 U$$726/A U$$764/B VGND VGND VPWR VPWR U$$726/X sky130_fd_sc_hd__xor2_1
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$737 U$$50/B1 U$$771/A2 U$$739/A1 U$$771/B2 VGND VGND VPWR VPWR U$$738/A sky130_fd_sc_hd__a22o_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$748 U$$748/A U$$774/B VGND VGND VPWR VPWR U$$748/X sky130_fd_sc_hd__xor2_1
XU$$759 U$$896/A1 U$$763/A2 U$$898/A1 U$$763/B2 VGND VGND VPWR VPWR U$$760/A sky130_fd_sc_hd__a22o_1
XFILLER_83_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_71_1 dadda_fa_3_71_1/A dadda_fa_3_71_1/B dadda_fa_3_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_0/CIN dadda_fa_4_71_2/A sky130_fd_sc_hd__fa_1
XFILLER_79_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_64_0 dadda_fa_3_64_0/A dadda_fa_3_64_0/B dadda_fa_3_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_0/B dadda_fa_4_64_1/CIN sky130_fd_sc_hd__fa_1
Xfanout1010 fanout1011/X VGND VGND VPWR VPWR U$$4458/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1021 U$$1189/B VGND VGND VPWR VPWR U$$1195/B sky130_fd_sc_hd__buf_6
Xfanout1032 U$$4315/B1 VGND VGND VPWR VPWR U$$479/B1 sky130_fd_sc_hd__buf_4
Xfanout1043 U$$4452/A1 VGND VGND VPWR VPWR U$$4315/A1 sky130_fd_sc_hd__buf_6
Xfanout1054 U$$66/A1 VGND VGND VPWR VPWR U$$64/B1 sky130_fd_sc_hd__buf_4
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1065 U$$612/A1 VGND VGND VPWR VPWR U$$747/B1 sky130_fd_sc_hd__buf_4
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1076 U$$4446/A1 VGND VGND VPWR VPWR U$$4309/A1 sky130_fd_sc_hd__buf_6
Xfanout1087 U$$3072/A1 VGND VGND VPWR VPWR U$$56/B1 sky130_fd_sc_hd__buf_4
XFILLER_48_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1098 input81/X VGND VGND VPWR VPWR U$$878/A1 sky130_fd_sc_hd__buf_6
XU$$2100 U$$2100/A U$$2130/B VGND VGND VPWR VPWR U$$2100/X sky130_fd_sc_hd__xor2_1
XFILLER_47_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2111 U$$878/A1 U$$2147/A2 U$$878/B1 U$$2147/B2 VGND VGND VPWR VPWR U$$2112/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_100_1 dadda_fa_4_100_1/A dadda_fa_4_100_1/B dadda_fa_4_100_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_101_0/B dadda_fa_5_100_1/B sky130_fd_sc_hd__fa_1
XFILLER_19_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2122 U$$2122/A U$$2130/B VGND VGND VPWR VPWR U$$2122/X sky130_fd_sc_hd__xor2_1
XU$$2133 U$$3775/B1 U$$2177/A2 U$$3642/A1 U$$2177/B2 VGND VGND VPWR VPWR U$$2134/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2144 U$$2144/A U$$2191/A VGND VGND VPWR VPWR U$$2144/X sky130_fd_sc_hd__xor2_1
XFILLER_35_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1410 U$$314/A1 U$$1452/A2 U$$42/A1 U$$1452/B2 VGND VGND VPWR VPWR U$$1411/A sky130_fd_sc_hd__a22o_1
XU$$2155 U$$3249/B1 U$$2181/A2 U$$4486/A1 U$$2181/B2 VGND VGND VPWR VPWR U$$2156/A
+ sky130_fd_sc_hd__a22o_1
XU$$1421 U$$1421/A U$$1427/B VGND VGND VPWR VPWR U$$1421/X sky130_fd_sc_hd__xor2_1
XU$$2166 U$$2166/A U$$2168/B VGND VGND VPWR VPWR U$$2166/X sky130_fd_sc_hd__xor2_1
XU$$1432 U$$884/A1 U$$1432/A2 U$$884/B1 U$$1432/B2 VGND VGND VPWR VPWR U$$1433/A sky130_fd_sc_hd__a22o_1
XU$$2177 U$$2860/B1 U$$2177/A2 U$$2862/B1 U$$2177/B2 VGND VGND VPWR VPWR U$$2178/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4463_1879 VGND VGND VPWR VPWR U$$4463_1879/HI U$$4463/B sky130_fd_sc_hd__conb_1
XU$$2188 U$$2188/A U$$2191/A VGND VGND VPWR VPWR U$$2188/X sky130_fd_sc_hd__xor2_1
XU$$1443 U$$1443/A U$$1449/B VGND VGND VPWR VPWR U$$1443/X sky130_fd_sc_hd__xor2_1
XU$$2199 U$$2199/A U$$2231/B VGND VGND VPWR VPWR U$$2199/X sky130_fd_sc_hd__xor2_1
XU$$1454 U$$82/B1 U$$1480/A2 U$$906/B1 U$$1480/B2 VGND VGND VPWR VPWR U$$1455/A sky130_fd_sc_hd__a22o_1
XU$$1465 U$$1465/A U$$1475/B VGND VGND VPWR VPWR U$$1465/X sky130_fd_sc_hd__xor2_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1476 U$$654/A1 U$$1480/A2 U$$654/B1 U$$1480/B2 VGND VGND VPWR VPWR U$$1477/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_7_121_0 dadda_fa_7_121_0/A dadda_fa_7_121_0/B dadda_fa_7_121_0/CIN VGND
+ VGND VPWR VPWR _418_/D _289_/D sky130_fd_sc_hd__fa_1
XU$$1487 U$$1487/A U$$1491/B VGND VGND VPWR VPWR U$$1487/X sky130_fd_sc_hd__xor2_1
XU$$1498 U$$539/A1 U$$1504/A2 U$$539/B1 U$$1504/B2 VGND VGND VPWR VPWR U$$1499/A sky130_fd_sc_hd__a22o_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_106_0_1934 VGND VGND VPWR VPWR dadda_fa_2_106_0/A dadda_fa_2_106_0_1934/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_31_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_86_1 dadda_fa_5_86_1/A dadda_fa_5_86_1/B dadda_fa_5_86_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_87_0/B dadda_fa_7_86_0/A sky130_fd_sc_hd__fa_2
XFILLER_7_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_79_0 dadda_fa_5_79_0/A dadda_fa_5_79_0/B dadda_fa_5_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_80_0/A dadda_fa_6_79_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_171_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_78_8 U$$4419/X input232/X dadda_fa_1_78_8/CIN VGND VGND VPWR VPWR dadda_fa_2_79_3/A
+ dadda_fa_3_78_0/A sky130_fd_sc_hd__fa_2
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$106 _402_/Q _274_/Q VGND VGND VPWR VPWR final_adder.U$$919/B1 final_adder.U$$148/A
+ sky130_fd_sc_hd__ha_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$117 _413_/Q _285_/Q VGND VGND VPWR VPWR final_adder.U$$139/B1 final_adder.U$$138/B
+ sky130_fd_sc_hd__ha_1
XFILLER_39_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$139 final_adder.U$$138/B final_adder.U$$909/B1 final_adder.U$$139/B1
+ VGND VGND VPWR VPWR final_adder.U$$139/X sky130_fd_sc_hd__a21o_1
XFILLER_39_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4080 U$$4080/A U$$4082/B VGND VGND VPWR VPWR U$$4080/X sky130_fd_sc_hd__xor2_1
XFILLER_26_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4091 U$$4226/B1 U$$4093/A2 U$$4093/A1 U$$4093/B2 VGND VGND VPWR VPWR U$$4092/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3390 U$$650/A1 U$$3390/A2 U$$650/B1 U$$3390/B2 VGND VGND VPWR VPWR U$$3391/A sky130_fd_sc_hd__a22o_1
XFILLER_13_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_81_0 dadda_fa_4_81_0/A dadda_fa_4_81_0/B dadda_fa_4_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_82_0/A dadda_fa_5_81_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_102_3 dadda_fa_3_102_3/A dadda_fa_3_102_3/B dadda_fa_3_102_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_103_1/B dadda_fa_4_102_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_70_0_1919 VGND VGND VPWR VPWR dadda_fa_0_70_0/A dadda_fa_0_70_0_1919/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_89_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput102 b[43] VGND VGND VPWR VPWR input102/X sky130_fd_sc_hd__buf_2
XFILLER_103_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput113 b[53] VGND VGND VPWR VPWR input113/X sky130_fd_sc_hd__clkbuf_1
Xinput124 b[63] VGND VGND VPWR VPWR input124/X sky130_fd_sc_hd__buf_4
XFILLER_131_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput135 c[105] VGND VGND VPWR VPWR input135/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput146 c[115] VGND VGND VPWR VPWR input146/X sky130_fd_sc_hd__clkbuf_4
Xinput157 c[125] VGND VGND VPWR VPWR input157/X sky130_fd_sc_hd__clkbuf_2
Xinput168 c[1] VGND VGND VPWR VPWR input168/X sky130_fd_sc_hd__clkbuf_4
Xfinal_adder.U$$640 final_adder.U$$656/B final_adder.U$$640/B VGND VGND VPWR VPWR
+ final_adder.U$$752/B sky130_fd_sc_hd__and2_1
Xinput179 c[2] VGND VGND VPWR VPWR input179/X sky130_fd_sc_hd__clkbuf_4
Xfinal_adder.U$$651 final_adder.U$$650/B final_adder.U$$547/X final_adder.U$$531/X
+ VGND VGND VPWR VPWR final_adder.U$$651/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$662 final_adder.U$$678/B final_adder.U$$662/B VGND VGND VPWR VPWR
+ final_adder.U$$774/B sky130_fd_sc_hd__and2_1
XU$$501 U$$88/B1 U$$501/A2 U$$503/A1 U$$501/B2 VGND VGND VPWR VPWR U$$502/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_109_0 dadda_fa_6_109_0/A dadda_fa_6_109_0/B dadda_fa_6_109_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_110_0/B dadda_fa_7_109_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$673 final_adder.U$$672/B final_adder.U$$569/X final_adder.U$$553/X
+ VGND VGND VPWR VPWR final_adder.U$$673/X sky130_fd_sc_hd__a21o_1
XFILLER_29_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$512 U$$512/A U$$522/B VGND VGND VPWR VPWR U$$512/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$684 final_adder.U$$700/B final_adder.U$$684/B VGND VGND VPWR VPWR
+ final_adder.U$$796/B sky130_fd_sc_hd__and2_1
XU$$523 U$$934/A1 U$$539/A2 U$$936/A1 U$$539/B2 VGND VGND VPWR VPWR U$$524/A sky130_fd_sc_hd__a22o_1
XFILLER_72_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$695 final_adder.U$$694/B final_adder.U$$591/X final_adder.U$$575/X
+ VGND VGND VPWR VPWR final_adder.U$$695/X sky130_fd_sc_hd__a21o_1
XU$$534 U$$534/A U$$536/B VGND VGND VPWR VPWR U$$534/X sky130_fd_sc_hd__xor2_1
XFILLER_17_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$545 U$$545/A1 U$$545/A2 U$$545/B1 U$$545/B2 VGND VGND VPWR VPWR U$$546/A sky130_fd_sc_hd__a22o_1
XU$$556 U$$965/B1 U$$610/A2 U$$10/A1 U$$610/B2 VGND VGND VPWR VPWR U$$557/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_29_3 dadda_fa_3_29_3/A dadda_fa_3_29_3/B dadda_fa_3_29_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_30_1/B dadda_fa_4_29_2/CIN sky130_fd_sc_hd__fa_1
XU$$567 U$$567/A U$$607/B VGND VGND VPWR VPWR U$$567/X sky130_fd_sc_hd__xor2_1
XU$$578 U$$30/A1 U$$610/A2 U$$32/A1 U$$610/B2 VGND VGND VPWR VPWR U$$579/A sky130_fd_sc_hd__a22o_1
XU$$589 U$$589/A U$$631/B VGND VGND VPWR VPWR U$$589/X sky130_fd_sc_hd__xor2_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_96_0 dadda_fa_6_96_0/A dadda_fa_6_96_0/B dadda_fa_6_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_97_0/B dadda_fa_7_96_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_32_5 U$$2066/X U$$2199/X VGND VGND VPWR VPWR dadda_fa_3_33_2/A dadda_fa_4_32_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_94_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_31_3 U$$1266/X U$$1399/X U$$1532/X VGND VGND VPWR VPWR dadda_fa_3_32_1/CIN
+ dadda_fa_3_31_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1240 U$$1240/A U$$1282/B VGND VGND VPWR VPWR U$$1240/X sky130_fd_sc_hd__xor2_1
XFILLER_22_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1251 U$$3030/B1 U$$1327/A2 U$$2897/A1 U$$1327/B2 VGND VGND VPWR VPWR U$$1252/A
+ sky130_fd_sc_hd__a22o_1
XU$$1262 U$$1262/A U$$1294/B VGND VGND VPWR VPWR U$$1262/X sky130_fd_sc_hd__xor2_1
XU$$1273 U$$314/A1 U$$1309/A2 U$$42/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1274/A sky130_fd_sc_hd__a22o_1
XU$$1284 U$$1284/A U$$1300/B VGND VGND VPWR VPWR U$$1284/X sky130_fd_sc_hd__xor2_1
XU$$1295 U$$62/A1 U$$1295/A2 U$$64/A1 U$$1295/B2 VGND VGND VPWR VPWR U$$1296/A sky130_fd_sc_hd__a22o_1
XFILLER_136_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_6 U$$3764/X U$$3897/X U$$4030/X VGND VGND VPWR VPWR dadda_fa_2_84_3/CIN
+ dadda_fa_3_83_0/A sky130_fd_sc_hd__fa_1
Xfanout803 U$$2745/X VGND VGND VPWR VPWR U$$2812/B2 sky130_fd_sc_hd__buf_4
Xfanout814 fanout820/X VGND VGND VPWR VPWR U$$2574/B2 sky130_fd_sc_hd__buf_6
Xfanout825 U$$2463/B2 VGND VGND VPWR VPWR U$$2415/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_131_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_76_5 U$$3484/X U$$3617/X U$$3750/X VGND VGND VPWR VPWR dadda_fa_2_77_2/A
+ dadda_fa_2_76_5/A sky130_fd_sc_hd__fa_1
Xfanout836 U$$2197/X VGND VGND VPWR VPWR U$$2320/B2 sky130_fd_sc_hd__buf_4
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout847 U$$2014/B2 VGND VGND VPWR VPWR U$$1980/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout858 U$$1915/B2 VGND VGND VPWR VPWR U$$1909/B2 sky130_fd_sc_hd__buf_6
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout869 U$$1760/B2 VGND VGND VPWR VPWR U$$1758/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_69_4 U$$4002/X U$$4135/X U$$4268/X VGND VGND VPWR VPWR dadda_fa_2_70_1/CIN
+ dadda_fa_2_69_4/CIN sky130_fd_sc_hd__fa_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_39_2 dadda_fa_4_39_2/A dadda_fa_4_39_2/B dadda_fa_4_39_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_40_0/CIN dadda_fa_5_39_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4485_1890 VGND VGND VPWR VPWR U$$4485_1890/HI U$$4485/B sky130_fd_sc_hd__conb_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_100_0 U$$4330/X U$$4463/X input130/X VGND VGND VPWR VPWR dadda_fa_4_101_0/B
+ dadda_fa_4_100_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_64_3 U$$1332/X U$$1465/X U$$1598/X VGND VGND VPWR VPWR dadda_fa_1_65_6/B
+ dadda_fa_1_64_8/B sky130_fd_sc_hd__fa_1
XFILLER_67_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_41_2 dadda_fa_3_41_2/A dadda_fa_3_41_2/B dadda_fa_3_41_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_1/A dadda_fa_4_41_2/B sky130_fd_sc_hd__fa_1
XFILLER_17_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$470 final_adder.U$$474/B final_adder.U$$470/B VGND VGND VPWR VPWR
+ final_adder.U$$594/B sky130_fd_sc_hd__and2_1
XFILLER_18_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$481 final_adder.U$$480/B final_adder.U$$359/X final_adder.U$$355/X
+ VGND VGND VPWR VPWR final_adder.U$$481/X sky130_fd_sc_hd__a21o_1
XU$$320 U$$868/A1 U$$352/A2 U$$868/B1 U$$352/B2 VGND VGND VPWR VPWR U$$321/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_34_1 dadda_fa_3_34_1/A dadda_fa_3_34_1/B dadda_fa_3_34_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_0/CIN dadda_fa_4_34_2/A sky130_fd_sc_hd__fa_1
XFILLER_123_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$492 final_adder.U$$496/B final_adder.U$$492/B VGND VGND VPWR VPWR
+ final_adder.U$$616/B sky130_fd_sc_hd__and2_1
XU$$331 U$$331/A U$$363/B VGND VGND VPWR VPWR U$$331/X sky130_fd_sc_hd__xor2_1
XU$$342 U$$479/A1 U$$346/A2 U$$481/A1 U$$346/B2 VGND VGND VPWR VPWR U$$343/A sky130_fd_sc_hd__a22o_1
XFILLER_18_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$353 U$$353/A U$$353/B VGND VGND VPWR VPWR U$$353/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_11_0 dadda_fa_6_11_0/A dadda_fa_6_11_0/B dadda_fa_6_11_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_12_0/B dadda_fa_7_11_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_27_0 U$$1125/X U$$1258/X U$$1391/X VGND VGND VPWR VPWR dadda_fa_4_28_0/B
+ dadda_fa_4_27_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_60_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$364 U$$90/A1 U$$406/A2 U$$92/A1 U$$406/B2 VGND VGND VPWR VPWR U$$365/A sky130_fd_sc_hd__a22o_1
XU$$375 U$$375/A U$$387/B VGND VGND VPWR VPWR U$$375/X sky130_fd_sc_hd__xor2_1
XU$$386 U$$521/B1 U$$386/A2 U$$386/B1 U$$386/B2 VGND VGND VPWR VPWR U$$387/A sky130_fd_sc_hd__a22o_1
XU$$397 U$$397/A U$$411/A VGND VGND VPWR VPWR U$$397/X sky130_fd_sc_hd__xor2_1
XFILLER_32_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_93_5 dadda_fa_2_93_5/A dadda_fa_2_93_5/B dadda_fa_2_93_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_94_2/A dadda_fa_4_93_0/A sky130_fd_sc_hd__fa_2
XFILLER_126_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_86_4 dadda_fa_2_86_4/A dadda_fa_2_86_4/B dadda_fa_2_86_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_87_1/CIN dadda_fa_3_86_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_79_3 dadda_fa_2_79_3/A dadda_fa_2_79_3/B dadda_fa_2_79_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_1/B dadda_fa_3_79_3/B sky130_fd_sc_hd__fa_1
XFILLER_67_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_49_1 dadda_fa_5_49_1/A dadda_fa_5_49_1/B dadda_fa_5_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_50_0/B dadda_fa_7_49_0/A sky130_fd_sc_hd__fa_1
XFILLER_79_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_102_2 U$$3403/X U$$3536/X U$$3669/X VGND VGND VPWR VPWR dadda_fa_3_103_2/CIN
+ dadda_fa_3_102_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_51_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1070 U$$1070/A U$$962/A VGND VGND VPWR VPWR U$$1070/X sky130_fd_sc_hd__xor2_1
XU$$1081 U$$120/B1 U$$1093/A2 U$$946/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1082/A sky130_fd_sc_hd__a22o_1
XFILLER_32_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1092 U$$1092/A U$$1094/B VGND VGND VPWR VPWR U$$1092/X sky130_fd_sc_hd__xor2_1
XFILLER_149_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_123_1 U$$4509/X input155/X dadda_fa_5_123_1/CIN VGND VGND VPWR VPWR dadda_fa_6_124_0/B
+ dadda_fa_7_123_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_116_0 dadda_fa_5_116_0/A dadda_fa_5_116_0/B dadda_fa_5_116_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_117_0/A dadda_fa_6_116_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_81_3 U$$2430/X U$$2563/X U$$2696/X VGND VGND VPWR VPWR dadda_fa_2_82_2/A
+ dadda_fa_2_81_4/CIN sky130_fd_sc_hd__fa_1
Xfanout600 U$$1915/A2 VGND VGND VPWR VPWR U$$1911/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout1609 input118/X VGND VGND VPWR VPWR U$$2862/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout611 U$$1648/X VGND VGND VPWR VPWR U$$1760/A2 sky130_fd_sc_hd__buf_6
Xfanout622 U$$259/A2 VGND VGND VPWR VPWR U$$219/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_74_2 U$$2549/X U$$2682/X U$$2815/X VGND VGND VPWR VPWR dadda_fa_2_75_1/A
+ dadda_fa_2_74_4/A sky130_fd_sc_hd__fa_1
XFILLER_77_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout633 U$$1480/A2 VGND VGND VPWR VPWR U$$1452/A2 sky130_fd_sc_hd__buf_6
Xfanout644 U$$1237/X VGND VGND VPWR VPWR U$$1353/A2 sky130_fd_sc_hd__buf_6
Xfanout655 U$$964/X VGND VGND VPWR VPWR U$$1075/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_4_51_1 dadda_fa_4_51_1/A dadda_fa_4_51_1/B dadda_fa_4_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_52_0/B dadda_fa_5_51_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_67_1 U$$2934/X U$$3067/X U$$3200/X VGND VGND VPWR VPWR dadda_fa_2_68_0/CIN
+ dadda_fa_2_67_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout666 U$$952/B2 VGND VGND VPWR VPWR U$$956/B2 sky130_fd_sc_hd__clkbuf_8
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout677 U$$676/B2 VGND VGND VPWR VPWR U$$636/B2 sky130_fd_sc_hd__buf_4
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout688 U$$4369/B2 VGND VGND VPWR VPWR U$$4349/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_44_0 dadda_fa_4_44_0/A dadda_fa_4_44_0/B dadda_fa_4_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_45_0/A dadda_fa_5_44_1/A sky130_fd_sc_hd__fa_1
XFILLER_59_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout699 U$$545/B2 VGND VGND VPWR VPWR U$$505/B2 sky130_fd_sc_hd__buf_4
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_410_ _416_/CLK _410_/D VGND VGND VPWR VPWR _410_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_341_ _342_/CLK _341_/D VGND VGND VPWR VPWR _341_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_272_ _402_/CLK _272_/D VGND VGND VPWR VPWR _272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_96_3 dadda_fa_3_96_3/A dadda_fa_3_96_3/B dadda_fa_3_96_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_1/B dadda_fa_4_96_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_154_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_89_2 dadda_fa_3_89_2/A dadda_fa_3_89_2/B dadda_fa_3_89_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_1/A dadda_fa_4_89_2/B sky130_fd_sc_hd__fa_1
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_59_0 dadda_fa_6_59_0/A dadda_fa_6_59_0/B dadda_fa_6_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_60_0/B dadda_fa_7_59_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_62_0 U$$131/X U$$264/X U$$397/X VGND VGND VPWR VPWR dadda_fa_1_63_5/B
+ dadda_fa_1_62_7/B sky130_fd_sc_hd__fa_1
XFILLER_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3901 U$$3901/A U$$3907/B VGND VGND VPWR VPWR U$$3901/X sky130_fd_sc_hd__xor2_1
XFILLER_37_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3912 U$$4049/A1 U$$3912/A2 U$$4462/A1 U$$3912/B2 VGND VGND VPWR VPWR U$$3913/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3923 U$$3923/A U$$3925/B VGND VGND VPWR VPWR U$$3923/X sky130_fd_sc_hd__xor2_1
XFILLER_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3934 U$$4482/A1 U$$3960/A2 U$$4484/A1 U$$3960/B2 VGND VGND VPWR VPWR U$$3935/A
+ sky130_fd_sc_hd__a22o_1
XU$$3945 U$$3945/A U$$3949/B VGND VGND VPWR VPWR U$$3945/X sky130_fd_sc_hd__xor2_1
XU$$3956 U$$4093/A1 U$$3970/A2 U$$4093/B1 U$$3970/B2 VGND VGND VPWR VPWR U$$3957/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3967 U$$3967/A U$$3972/A VGND VGND VPWR VPWR U$$3967/X sky130_fd_sc_hd__xor2_1
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3978 U$$3976/B U$$3973/A input54/X U$$3973/Y VGND VGND VPWR VPWR U$$3978/X sky130_fd_sc_hd__a22o_2
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3989 U$$4400/A1 U$$4025/A2 U$$4400/B1 U$$4025/B2 VGND VGND VPWR VPWR U$$3990/A
+ sky130_fd_sc_hd__a22o_1
XU$$150 U$$150/A U$$180/B VGND VGND VPWR VPWR U$$150/X sky130_fd_sc_hd__xor2_1
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$161 U$$24/A1 U$$213/A2 U$$26/A1 U$$213/B2 VGND VGND VPWR VPWR U$$162/A sky130_fd_sc_hd__a22o_1
XU$$172 U$$172/A U$$210/B VGND VGND VPWR VPWR U$$172/X sky130_fd_sc_hd__xor2_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$183 U$$183/A1 U$$219/A2 U$$48/A1 U$$219/B2 VGND VGND VPWR VPWR U$$184/A sky130_fd_sc_hd__a22o_1
XU$$194 U$$194/A U$$230/B VGND VGND VPWR VPWR U$$194/X sky130_fd_sc_hd__xor2_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_91_2 U$$3913/X U$$4046/X U$$4179/X VGND VGND VPWR VPWR dadda_fa_3_92_1/A
+ dadda_fa_3_91_3/A sky130_fd_sc_hd__fa_1
XFILLER_160_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_84_1 U$$4431/X input239/X dadda_fa_2_84_1/CIN VGND VGND VPWR VPWR dadda_fa_3_85_0/CIN
+ dadda_fa_3_84_2/CIN sky130_fd_sc_hd__fa_1
Xoutput258 output258/A VGND VGND VPWR VPWR o[100] sky130_fd_sc_hd__buf_2
Xoutput269 output269/A VGND VGND VPWR VPWR o[110] sky130_fd_sc_hd__buf_2
Xdadda_fa_5_61_0 dadda_fa_5_61_0/A dadda_fa_5_61_0/B dadda_fa_5_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_62_0/A dadda_fa_6_61_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_2_77_0 dadda_fa_2_77_0/A dadda_fa_2_77_0/B dadda_fa_2_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_0/B dadda_fa_3_77_2/B sky130_fd_sc_hd__fa_1
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_60_8 dadda_fa_1_60_8/A dadda_fa_1_60_8/B dadda_fa_1_60_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_61_3/A dadda_fa_3_60_0/A sky130_fd_sc_hd__fa_2
XFILLER_67_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_53_7 U$$3172/X U$$3305/X U$$3438/X VGND VGND VPWR VPWR dadda_fa_2_54_2/CIN
+ dadda_fa_2_53_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_99_1 dadda_fa_4_99_1/A dadda_fa_4_99_1/B dadda_fa_4_99_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_100_0/B dadda_fa_5_99_1/B sky130_fd_sc_hd__fa_1
XFILLER_136_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_76_0 dadda_fa_7_76_0/A dadda_fa_7_76_0/B dadda_fa_7_76_0/CIN VGND VGND
+ VPWR VPWR _373_/D _244_/D sky130_fd_sc_hd__fa_1
XFILLER_118_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1406 U$$2745/A2 VGND VGND VPWR VPWR U$$2678/B sky130_fd_sc_hd__buf_6
Xfanout1417 fanout1419/X VGND VGND VPWR VPWR U$$2591/B sky130_fd_sc_hd__buf_8
Xfanout1428 input3/X VGND VGND VPWR VPWR U$$821/A sky130_fd_sc_hd__buf_8
Xfanout430 U$$505/A2 VGND VGND VPWR VPWR U$$479/A2 sky130_fd_sc_hd__clkbuf_2
Xfanout441 U$$102/A2 VGND VGND VPWR VPWR U$$96/A2 sky130_fd_sc_hd__buf_4
Xfanout1439 U$$2269/B VGND VGND VPWR VPWR U$$2231/B sky130_fd_sc_hd__buf_6
XFILLER_87_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout452 U$$4043/A2 VGND VGND VPWR VPWR U$$4045/A2 sky130_fd_sc_hd__buf_4
XFILLER_59_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout463 U$$3966/A2 VGND VGND VPWR VPWR U$$3970/A2 sky130_fd_sc_hd__buf_4
XFILLER_24_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout474 U$$3833/A2 VGND VGND VPWR VPWR U$$3825/A2 sky130_fd_sc_hd__buf_4
Xfanout485 U$$3511/A2 VGND VGND VPWR VPWR U$$3505/A2 sky130_fd_sc_hd__buf_4
XFILLER_74_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout496 U$$3292/X VGND VGND VPWR VPWR U$$3378/A2 sky130_fd_sc_hd__clkbuf_4
XU$$3208 U$$3208/A U$$3208/B VGND VGND VPWR VPWR U$$3208/X sky130_fd_sc_hd__xor2_1
XFILLER_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3219 U$$4315/A1 U$$3283/A2 U$$4454/A1 U$$3283/B2 VGND VGND VPWR VPWR U$$3220/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2507 U$$2507/A U$$2545/B VGND VGND VPWR VPWR U$$2507/X sky130_fd_sc_hd__xor2_1
XU$$2518 U$$735/B1 U$$2540/A2 U$$602/A1 U$$2540/B2 VGND VGND VPWR VPWR U$$2519/A sky130_fd_sc_hd__a22o_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2529 U$$2529/A U$$2529/B VGND VGND VPWR VPWR U$$2529/X sky130_fd_sc_hd__xor2_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1806 U$$1806/A U$$1836/B VGND VGND VPWR VPWR U$$1806/X sky130_fd_sc_hd__xor2_1
XU$$1817 U$$3322/B1 U$$1831/A2 U$$721/B1 U$$1831/B2 VGND VGND VPWR VPWR U$$1818/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1828 U$$1828/A U$$1828/B VGND VGND VPWR VPWR U$$1828/X sky130_fd_sc_hd__xor2_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1839 U$$880/A1 U$$1881/A2 U$$882/A1 U$$1881/B2 VGND VGND VPWR VPWR U$$1840/A sky130_fd_sc_hd__a22o_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_324_ _344_/CLK _324_/D VGND VGND VPWR VPWR _324_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_255_ _384_/CLK _255_/D VGND VGND VPWR VPWR _255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_186_ _321_/CLK _186_/D VGND VGND VPWR VPWR _186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_94_0 dadda_fa_3_94_0/A dadda_fa_3_94_0/B dadda_fa_3_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_0/B dadda_fa_4_94_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4410 U$$4410/A1 U$$4388/X U$$4412/A1 U$$4458/B2 VGND VGND VPWR VPWR U$$4411/A
+ sky130_fd_sc_hd__a22o_1
XU$$4421 U$$4421/A U$$4421/B VGND VGND VPWR VPWR U$$4421/X sky130_fd_sc_hd__xor2_1
XFILLER_93_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_56_5 dadda_fa_2_56_5/A dadda_fa_2_56_5/B dadda_fa_2_56_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_2/A dadda_fa_4_56_0/A sky130_fd_sc_hd__fa_1
XU$$4432 U$$4432/A1 U$$4388/X U$$4434/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4433/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4443 U$$4443/A U$$4443/B VGND VGND VPWR VPWR U$$4443/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_49_4 dadda_fa_2_49_4/A dadda_fa_2_49_4/B dadda_fa_2_49_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_1/CIN dadda_fa_3_49_3/CIN sky130_fd_sc_hd__fa_1
XU$$4454 U$$4454/A1 U$$4388/X U$$4456/A1 U$$4458/B2 VGND VGND VPWR VPWR U$$4455/A
+ sky130_fd_sc_hd__a22o_1
XU$$3720 U$$3720/A U$$3734/B VGND VGND VPWR VPWR U$$3720/X sky130_fd_sc_hd__xor2_1
XU$$4465 U$$4465/A U$$4465/B VGND VGND VPWR VPWR U$$4465/X sky130_fd_sc_hd__xor2_1
XU$$3731 U$$854/A1 U$$3757/A2 U$$3870/A1 U$$3757/B2 VGND VGND VPWR VPWR U$$3732/A
+ sky130_fd_sc_hd__a22o_1
XU$$4476 U$$4476/A1 U$$4388/X U$$4478/A1 U$$4488/B2 VGND VGND VPWR VPWR U$$4477/A
+ sky130_fd_sc_hd__a22o_1
XU$$3742 U$$3742/A U$$3790/B VGND VGND VPWR VPWR U$$3742/X sky130_fd_sc_hd__xor2_1
XU$$4487 U$$4487/A U$$4487/B VGND VGND VPWR VPWR U$$4487/X sky130_fd_sc_hd__xor2_1
XU$$3753 U$$4162/B1 U$$3773/A2 U$$4027/B1 U$$3773/B2 VGND VGND VPWR VPWR U$$3754/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4498 U$$4498/A1 U$$4388/X U$$4500/A1 U$$4506/B2 VGND VGND VPWR VPWR U$$4499/A
+ sky130_fd_sc_hd__a22o_1
XU$$3764 U$$3764/A U$$3774/B VGND VGND VPWR VPWR U$$3764/X sky130_fd_sc_hd__xor2_1
XFILLER_46_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3775 U$$3775/A1 U$$3777/A2 U$$3775/B1 U$$3777/B2 VGND VGND VPWR VPWR U$$3776/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3786 U$$3786/A U$$3816/B VGND VGND VPWR VPWR U$$3786/X sky130_fd_sc_hd__xor2_1
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3797 U$$4345/A1 U$$3825/A2 U$$4484/A1 U$$3825/B2 VGND VGND VPWR VPWR U$$3798/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_978 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_45_5 U$$2092/X U$$2225/X VGND VGND VPWR VPWR dadda_fa_2_46_3/CIN dadda_fa_3_45_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_51_4 U$$1705/X U$$1838/X U$$1971/X VGND VGND VPWR VPWR dadda_fa_2_52_1/CIN
+ dadda_fa_2_51_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$908 U$$908/A1 U$$910/A2 U$$910/A1 U$$910/B2 VGND VGND VPWR VPWR U$$909/A sky130_fd_sc_hd__a22o_1
XU$$919 U$$919/A U$$958/A VGND VGND VPWR VPWR U$$919/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_44_3 U$$1292/X U$$1425/X U$$1558/X VGND VGND VPWR VPWR dadda_fa_2_45_3/B
+ dadda_fa_2_44_5/B sky130_fd_sc_hd__fa_1
XFILLER_141_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_21_2 dadda_fa_4_21_2/A dadda_fa_4_21_2/B dadda_ha_3_21_3/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_22_0/CIN dadda_fa_5_21_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_14_1 U$$700/X U$$833/X U$$966/X VGND VGND VPWR VPWR dadda_fa_5_15_0/B
+ dadda_fa_5_14_1/B sky130_fd_sc_hd__fa_1
XFILLER_169_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_886 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1203 U$$854/B1 VGND VGND VPWR VPWR U$$856/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1214 U$$3181/B1 VGND VGND VPWR VPWR U$$443/A1 sky130_fd_sc_hd__buf_4
XFILLER_120_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1225 input67/X VGND VGND VPWR VPWR U$$4414/A1 sky130_fd_sc_hd__buf_6
Xfanout1236 U$$3981/A1 VGND VGND VPWR VPWR U$$4392/A1 sky130_fd_sc_hd__buf_4
Xfanout1247 U$$639/B VGND VGND VPWR VPWR U$$607/B sky130_fd_sc_hd__buf_6
Xfanout1258 U$$522/B VGND VGND VPWR VPWR U$$506/B sky130_fd_sc_hd__buf_6
Xdadda_fa_3_59_3 dadda_fa_3_59_3/A dadda_fa_3_59_3/B dadda_fa_3_59_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_1/B dadda_fa_4_59_2/CIN sky130_fd_sc_hd__fa_1
Xfanout1269 input60/X VGND VGND VPWR VPWR U$$4322/B sky130_fd_sc_hd__buf_6
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3005 U$$3825/B1 U$$3005/A2 U$$3692/A1 U$$3005/B2 VGND VGND VPWR VPWR U$$3006/A
+ sky130_fd_sc_hd__a22o_1
XU$$3016 U$$3107/B VGND VGND VPWR VPWR U$$3016/Y sky130_fd_sc_hd__inv_1
XU$$3027 U$$3027/A U$$3061/B VGND VGND VPWR VPWR U$$3027/X sky130_fd_sc_hd__xor2_1
XFILLER_47_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3038 U$$3447/B1 U$$3122/A2 U$$3314/A1 U$$3122/B2 VGND VGND VPWR VPWR U$$3039/A
+ sky130_fd_sc_hd__a22o_1
XU$$2304 U$$2576/B1 U$$2310/A2 U$$388/A1 U$$2310/B2 VGND VGND VPWR VPWR U$$2305/A
+ sky130_fd_sc_hd__a22o_1
XU$$3049 U$$3049/A U$$3077/B VGND VGND VPWR VPWR U$$3049/X sky130_fd_sc_hd__xor2_1
XFILLER_46_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2315 U$$2315/A U$$2328/A VGND VGND VPWR VPWR U$$2315/X sky130_fd_sc_hd__xor2_1
XU$$2326 U$$956/A1 U$$2326/A2 U$$2326/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2327/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2337 U$$967/A1 U$$2415/A2 U$$969/A1 U$$2415/B2 VGND VGND VPWR VPWR U$$2338/A sky130_fd_sc_hd__a22o_1
XU$$1603 U$$2973/A1 U$$1635/A2 U$$2973/B1 U$$1635/B2 VGND VGND VPWR VPWR U$$1604/A
+ sky130_fd_sc_hd__a22o_1
XU$$2348 U$$2348/A U$$2402/B VGND VGND VPWR VPWR U$$2348/X sky130_fd_sc_hd__xor2_1
XFILLER_61_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1614 U$$1614/A U$$1626/B VGND VGND VPWR VPWR U$$1614/X sky130_fd_sc_hd__xor2_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2359 U$$2631/B1 U$$2395/A2 U$$989/B1 U$$2395/B2 VGND VGND VPWR VPWR U$$2360/A
+ sky130_fd_sc_hd__a22o_1
XU$$1625 U$$253/B1 U$$1625/A2 U$$120/A1 U$$1625/B2 VGND VGND VPWR VPWR U$$1626/A sky130_fd_sc_hd__a22o_1
XU$$1636 U$$1636/A U$$1644/A VGND VGND VPWR VPWR U$$1636/X sky130_fd_sc_hd__xor2_1
XU$$1647 U$$1777/B U$$1647/B VGND VGND VPWR VPWR U$$1647/X sky130_fd_sc_hd__and2_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1658 U$$2754/A1 U$$1696/A2 U$$2891/B1 U$$1696/B2 VGND VGND VPWR VPWR U$$1659/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1669 U$$1669/A U$$1703/B VGND VGND VPWR VPWR U$$1669/X sky130_fd_sc_hd__xor2_1
XFILLER_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_307_ _321_/CLK _307_/D VGND VGND VPWR VPWR _307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_238_ _367_/CLK _238_/D VGND VGND VPWR VPWR _238_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_112_0_1937 VGND VGND VPWR VPWR dadda_fa_3_112_0/A dadda_fa_3_112_0_1937/LO
+ sky130_fd_sc_hd__conb_1
X_169_ _319_/CLK _169_/D VGND VGND VPWR VPWR _169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_61_3 dadda_fa_2_61_3/A dadda_fa_2_61_3/B dadda_fa_2_61_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_1/B dadda_fa_3_61_3/B sky130_fd_sc_hd__fa_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_54_2 dadda_fa_2_54_2/A dadda_fa_2_54_2/B dadda_fa_2_54_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_1/A dadda_fa_3_54_3/A sky130_fd_sc_hd__fa_1
Xfanout1770 input101/X VGND VGND VPWR VPWR U$$914/A1 sky130_fd_sc_hd__buf_4
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_31_1 dadda_fa_5_31_1/A dadda_fa_5_31_1/B dadda_fa_5_31_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_32_0/B dadda_fa_7_31_0/A sky130_fd_sc_hd__fa_1
XFILLER_66_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4240 U$$4375/B1 U$$4240/A2 U$$4240/B1 U$$4240/B2 VGND VGND VPWR VPWR U$$4241/A
+ sky130_fd_sc_hd__a22o_1
XU$$4251 U$$4249/Y input59/X U$$4247/A U$$4250/X U$$4247/Y VGND VGND VPWR VPWR U$$4251/X
+ sky130_fd_sc_hd__a32o_1
XU$$4262 U$$4262/A U$$4292/B VGND VGND VPWR VPWR U$$4262/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_47_1 U$$3160/X input198/X dadda_fa_2_47_1/CIN VGND VGND VPWR VPWR dadda_fa_3_48_0/CIN
+ dadda_fa_3_47_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4273 U$$4410/A1 U$$4325/A2 U$$4412/A1 U$$4325/B2 VGND VGND VPWR VPWR U$$4274/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_24_0 dadda_fa_5_24_0/A dadda_fa_5_24_0/B dadda_fa_5_24_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_25_0/A dadda_fa_6_24_0/CIN sky130_fd_sc_hd__fa_1
XU$$4284 U$$4284/A U$$4368/B VGND VGND VPWR VPWR U$$4284/X sky130_fd_sc_hd__xor2_1
XU$$4295 U$$4432/A1 U$$4295/A2 U$$4295/B1 U$$4295/B2 VGND VGND VPWR VPWR U$$4296/A
+ sky130_fd_sc_hd__a22o_1
XU$$3550 U$$3550/A U$$3558/B VGND VGND VPWR VPWR U$$3550/X sky130_fd_sc_hd__xor2_1
XFILLER_25_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3561 U$$3561/A VGND VGND VPWR VPWR U$$3561/Y sky130_fd_sc_hd__inv_1
XU$$3572 U$$3846/A1 U$$3658/A2 U$$3846/B1 U$$3658/B2 VGND VGND VPWR VPWR U$$3573/A
+ sky130_fd_sc_hd__a22o_1
XU$$3583 U$$3583/A U$$3607/B VGND VGND VPWR VPWR U$$3583/X sky130_fd_sc_hd__xor2_1
XU$$3594 U$$854/A1 U$$3604/A2 U$$3870/A1 U$$3604/B2 VGND VGND VPWR VPWR U$$3595/A
+ sky130_fd_sc_hd__a22o_1
XU$$2860 U$$2860/A1 U$$2872/A2 U$$2860/B1 U$$2872/B2 VGND VGND VPWR VPWR U$$2861/A
+ sky130_fd_sc_hd__a22o_1
XU$$2871 U$$2871/A U$$2871/B VGND VGND VPWR VPWR U$$2871/X sky130_fd_sc_hd__xor2_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2882 U$$2880/B U$$2877/A input37/X U$$2877/Y VGND VGND VPWR VPWR U$$2882/X sky130_fd_sc_hd__a22o_4
XU$$2893 U$$3030/A1 U$$2929/A2 U$$3030/B1 U$$2929/B2 VGND VGND VPWR VPWR U$$2894/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_69_2 dadda_fa_4_69_2/A dadda_fa_4_69_2/B dadda_fa_4_69_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_70_0/CIN dadda_fa_5_69_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$800 final_adder.U$$800/A final_adder.U$$800/B VGND VGND VPWR VPWR
+ final_adder.U$$800/X sky130_fd_sc_hd__and2_1
XFILLER_102_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_36_1 U$$478/X U$$611/X VGND VGND VPWR VPWR dadda_fa_2_37_5/B dadda_fa_3_36_0/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$811 final_adder.U$$778/A final_adder.U$$731/X final_adder.U$$699/X
+ VGND VGND VPWR VPWR final_adder.U$$811/X sky130_fd_sc_hd__a21o_1
XFILLER_57_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_39_0 dadda_fa_7_39_0/A dadda_fa_7_39_0/B dadda_fa_7_39_0/CIN VGND VGND
+ VPWR VPWR _336_/D _207_/D sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$833 final_adder.U$$800/A final_adder.U$$255/X final_adder.U$$721/X
+ VGND VGND VPWR VPWR final_adder.U$$833/X sky130_fd_sc_hd__a21o_1
XFILLER_21_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$855 final_adder.U$$758/X final_adder.U$$823/X final_adder.U$$759/X
+ VGND VGND VPWR VPWR final_adder.U$$855/X sky130_fd_sc_hd__a21o_1
XU$$705 U$$840/B1 U$$771/A2 U$$707/A1 U$$771/B2 VGND VGND VPWR VPWR U$$706/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$877 final_adder.U$$780/X final_adder.U$$733/X final_adder.U$$781/X
+ VGND VGND VPWR VPWR final_adder.U$$877/X sky130_fd_sc_hd__a21o_1
XU$$716 U$$716/A U$$774/B VGND VGND VPWR VPWR U$$716/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_42_0 U$$91/X U$$224/X U$$357/X VGND VGND VPWR VPWR dadda_fa_2_43_3/A dadda_fa_2_42_4/CIN
+ sky130_fd_sc_hd__fa_1
XU$$727 U$$864/A1 U$$763/A2 U$$864/B1 U$$763/B2 VGND VGND VPWR VPWR U$$728/A sky130_fd_sc_hd__a22o_1
XU$$738 U$$738/A U$$774/B VGND VGND VPWR VPWR U$$738/X sky130_fd_sc_hd__xor2_1
XU$$4449_1872 VGND VGND VPWR VPWR U$$4449_1872/HI U$$4449/B sky130_fd_sc_hd__conb_1
XFILLER_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$899 final_adder.U$$899/A1 final_adder.U$$837/X final_adder.U$$899/B1
+ VGND VGND VPWR VPWR final_adder.U$$899/X sky130_fd_sc_hd__a21o_1
XFILLER_72_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$749 U$$884/B1 U$$769/A2 U$$749/B1 U$$769/B2 VGND VGND VPWR VPWR U$$750/A sky130_fd_sc_hd__a22o_1
XFILLER_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_71_2 dadda_fa_3_71_2/A dadda_fa_3_71_2/B dadda_fa_3_71_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_1/A dadda_fa_4_71_2/B sky130_fd_sc_hd__fa_1
Xfanout1000 fanout999/A VGND VGND VPWR VPWR U$$4049/A1 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_3_64_1 dadda_fa_3_64_1/A dadda_fa_3_64_1/B dadda_fa_3_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_0/CIN dadda_fa_4_64_2/A sky130_fd_sc_hd__fa_1
Xfanout1011 input91/X VGND VGND VPWR VPWR fanout1011/X sky130_fd_sc_hd__buf_6
XFILLER_126_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1022 U$$1189/B VGND VGND VPWR VPWR U$$1233/A sky130_fd_sc_hd__buf_4
XFILLER_0_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1033 U$$4315/B1 VGND VGND VPWR VPWR U$$3630/B1 sky130_fd_sc_hd__buf_4
XFILLER_121_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_41_0 dadda_fa_6_41_0/A dadda_fa_6_41_0/B dadda_fa_6_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_42_0/B dadda_fa_7_41_0/CIN sky130_fd_sc_hd__fa_1
Xfanout1044 input88/X VGND VGND VPWR VPWR U$$4452/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout1055 U$$3080/A1 VGND VGND VPWR VPWR U$$66/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_57_0 dadda_fa_3_57_0/A dadda_fa_3_57_0/B dadda_fa_3_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_0/B dadda_fa_4_57_1/CIN sky130_fd_sc_hd__fa_1
Xfanout1066 input85/X VGND VGND VPWR VPWR U$$612/A1 sky130_fd_sc_hd__buf_6
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1077 input84/X VGND VGND VPWR VPWR U$$4446/A1 sky130_fd_sc_hd__buf_4
Xfanout1088 input82/X VGND VGND VPWR VPWR U$$3072/A1 sky130_fd_sc_hd__buf_4
Xfanout1099 U$$3618/A1 VGND VGND VPWR VPWR U$$4027/B1 sky130_fd_sc_hd__buf_6
XFILLER_48_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2101 U$$183/A1 U$$2107/A2 U$$870/A1 U$$2107/B2 VGND VGND VPWR VPWR U$$2102/A sky130_fd_sc_hd__a22o_1
XU$$2112 U$$2112/A U$$2148/B VGND VGND VPWR VPWR U$$2112/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_100_2 dadda_fa_4_100_2/A dadda_fa_4_100_2/B dadda_fa_4_100_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_101_0/CIN dadda_fa_5_100_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2123 U$$68/A1 U$$2139/A2 U$$70/A1 U$$2139/B2 VGND VGND VPWR VPWR U$$2124/A sky130_fd_sc_hd__a22o_1
XU$$2134 U$$2134/A U$$2168/B VGND VGND VPWR VPWR U$$2134/X sky130_fd_sc_hd__xor2_1
XFILLER_62_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1400 U$$2631/B1 U$$1414/A2 U$$852/B1 U$$1414/B2 VGND VGND VPWR VPWR U$$1401/A
+ sky130_fd_sc_hd__a22o_1
XU$$2145 U$$773/B1 U$$2147/A2 U$$640/A1 U$$2147/B2 VGND VGND VPWR VPWR U$$2146/A sky130_fd_sc_hd__a22o_1
XU$$1411 U$$1411/A U$$1449/B VGND VGND VPWR VPWR U$$1411/X sky130_fd_sc_hd__xor2_1
XU$$2156 U$$2156/A U$$2191/A VGND VGND VPWR VPWR U$$2156/X sky130_fd_sc_hd__xor2_1
XU$$1422 U$$598/B1 U$$1426/A2 U$$465/A1 U$$1426/B2 VGND VGND VPWR VPWR U$$1423/A sky130_fd_sc_hd__a22o_1
XU$$2167 U$$2576/B1 U$$2181/A2 U$$388/A1 U$$2181/B2 VGND VGND VPWR VPWR U$$2168/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1433 U$$1433/A U$$1433/B VGND VGND VPWR VPWR U$$1433/X sky130_fd_sc_hd__xor2_1
XU$$2178 U$$2178/A U$$2192/A VGND VGND VPWR VPWR U$$2178/X sky130_fd_sc_hd__xor2_1
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2189 U$$3833/A1 U$$2189/A2 U$$2189/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2190/A
+ sky130_fd_sc_hd__a22o_1
XU$$1444 U$$2814/A1 U$$1452/A2 U$$76/A1 U$$1452/B2 VGND VGND VPWR VPWR U$$1445/A sky130_fd_sc_hd__a22o_1
XFILLER_71_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1455 U$$1455/A U$$1455/B VGND VGND VPWR VPWR U$$1455/X sky130_fd_sc_hd__xor2_1
XU$$1466 U$$2973/A1 U$$1502/A2 U$$2973/B1 U$$1502/B2 VGND VGND VPWR VPWR U$$1467/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1477 U$$1477/A U$$1491/B VGND VGND VPWR VPWR U$$1477/X sky130_fd_sc_hd__xor2_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1488 U$$4365/A1 U$$1502/A2 U$$4365/B1 U$$1502/B2 VGND VGND VPWR VPWR U$$1489/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1499 U$$1499/A U$$1507/A VGND VGND VPWR VPWR U$$1499/X sky130_fd_sc_hd__xor2_1
XFILLER_124_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_114_0 dadda_fa_7_114_0/A dadda_fa_7_114_0/B dadda_fa_7_114_0/CIN VGND
+ VGND VPWR VPWR _411_/D _282_/D sky130_fd_sc_hd__fa_1
XFILLER_128_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_79_1 dadda_fa_5_79_1/A dadda_fa_5_79_1/B dadda_fa_5_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_80_0/B dadda_fa_7_79_0/A sky130_fd_sc_hd__fa_2
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$107 _403_/Q _275_/Q VGND VGND VPWR VPWR final_adder.U$$149/B1 final_adder.U$$148/B
+ sky130_fd_sc_hd__ha_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$118 _414_/Q _286_/Q VGND VGND VPWR VPWR final_adder.U$$907/B1 final_adder.U$$136/A
+ sky130_fd_sc_hd__ha_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4070 U$$4070/A U$$4082/B VGND VGND VPWR VPWR U$$4070/X sky130_fd_sc_hd__xor2_1
XFILLER_66_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4081 U$$4081/A1 U$$4081/A2 U$$4081/B1 U$$4081/B2 VGND VGND VPWR VPWR U$$4082/A
+ sky130_fd_sc_hd__a22o_1
XU$$4092 U$$4092/A U$$4094/B VGND VGND VPWR VPWR U$$4092/X sky130_fd_sc_hd__xor2_1
XFILLER_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3380 U$$3515/B1 U$$3422/A2 U$$3382/A1 U$$3422/B2 VGND VGND VPWR VPWR U$$3381/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3391 U$$3391/A U$$3391/B VGND VGND VPWR VPWR U$$3391/X sky130_fd_sc_hd__xor2_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2690 U$$2690/A U$$2740/A VGND VGND VPWR VPWR U$$2690/X sky130_fd_sc_hd__xor2_1
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4479_1887 VGND VGND VPWR VPWR U$$4479_1887/HI U$$4479/B sky130_fd_sc_hd__conb_1
XFILLER_147_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_81_1 dadda_fa_4_81_1/A dadda_fa_4_81_1/B dadda_fa_4_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_82_0/B dadda_fa_5_81_1/B sky130_fd_sc_hd__fa_1
XFILLER_89_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_74_0 dadda_fa_4_74_0/A dadda_fa_4_74_0/B dadda_fa_4_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_75_0/A dadda_fa_5_74_1/A sky130_fd_sc_hd__fa_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput103 b[44] VGND VGND VPWR VPWR input103/X sky130_fd_sc_hd__buf_2
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput114 b[54] VGND VGND VPWR VPWR input114/X sky130_fd_sc_hd__buf_4
XFILLER_49_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput125 b[6] VGND VGND VPWR VPWR input125/X sky130_fd_sc_hd__buf_2
Xinput136 c[106] VGND VGND VPWR VPWR input136/X sky130_fd_sc_hd__clkbuf_4
Xinput147 c[116] VGND VGND VPWR VPWR input147/X sky130_fd_sc_hd__clkbuf_4
Xinput158 c[126] VGND VGND VPWR VPWR input158/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput169 c[20] VGND VGND VPWR VPWR input169/X sky130_fd_sc_hd__clkbuf_4
Xfinal_adder.U$$630 final_adder.U$$646/B final_adder.U$$630/B VGND VGND VPWR VPWR
+ final_adder.U$$742/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$641 final_adder.U$$640/B final_adder.U$$537/X final_adder.U$$521/X
+ VGND VGND VPWR VPWR final_adder.U$$641/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$652 final_adder.U$$668/B final_adder.U$$652/B VGND VGND VPWR VPWR
+ final_adder.U$$764/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$663 final_adder.U$$662/B final_adder.U$$559/X final_adder.U$$543/X
+ VGND VGND VPWR VPWR final_adder.U$$663/X sky130_fd_sc_hd__a21o_1
XU$$502 U$$502/A U$$504/B VGND VGND VPWR VPWR U$$502/X sky130_fd_sc_hd__xor2_1
XFILLER_91_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$674 final_adder.U$$690/B final_adder.U$$674/B VGND VGND VPWR VPWR
+ final_adder.U$$786/B sky130_fd_sc_hd__and2_1
XU$$513 U$$650/A1 U$$415/X U$$650/B1 U$$416/X VGND VGND VPWR VPWR U$$514/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$685 final_adder.U$$684/B final_adder.U$$581/X final_adder.U$$565/X
+ VGND VGND VPWR VPWR final_adder.U$$685/X sky130_fd_sc_hd__a21o_1
XU$$524 U$$524/A U$$536/B VGND VGND VPWR VPWR U$$524/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$696 final_adder.U$$712/B final_adder.U$$696/B VGND VGND VPWR VPWR
+ final_adder.U$$776/A sky130_fd_sc_hd__and2_1
XU$$535 U$$672/A1 U$$539/A2 U$$672/B1 U$$539/B2 VGND VGND VPWR VPWR U$$536/A sky130_fd_sc_hd__a22o_1
XU$$546 U$$546/A U$$547/A VGND VGND VPWR VPWR U$$546/X sky130_fd_sc_hd__xor2_1
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$557 U$$557/A U$$607/B VGND VGND VPWR VPWR U$$557/X sky130_fd_sc_hd__xor2_1
XFILLER_60_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$568 U$$840/B1 U$$638/A2 U$$707/A1 U$$638/B2 VGND VGND VPWR VPWR U$$569/A sky130_fd_sc_hd__a22o_1
XU$$579 U$$579/A U$$607/B VGND VGND VPWR VPWR U$$579/X sky130_fd_sc_hd__xor2_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_89_0 dadda_fa_6_89_0/A dadda_fa_6_89_0/B dadda_fa_6_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_90_0/B dadda_fa_7_89_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_172_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1230 U$$406/B1 U$$1230/A2 U$$1230/B1 U$$1230/B2 VGND VGND VPWR VPWR U$$1231/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1241 U$$967/A1 U$$1311/A2 U$$969/A1 U$$1311/B2 VGND VGND VPWR VPWR U$$1242/A sky130_fd_sc_hd__a22o_1
XU$$1252 U$$1252/A U$$1294/B VGND VGND VPWR VPWR U$$1252/X sky130_fd_sc_hd__xor2_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1263 U$$989/A1 U$$1327/A2 U$$991/A1 U$$1327/B2 VGND VGND VPWR VPWR U$$1264/A sky130_fd_sc_hd__a22o_1
XU$$1274 U$$1274/A U$$1278/B VGND VGND VPWR VPWR U$$1274/X sky130_fd_sc_hd__xor2_1
XU$$1285 U$$52/A1 U$$1327/A2 U$$54/A1 U$$1327/B2 VGND VGND VPWR VPWR U$$1286/A sky130_fd_sc_hd__a22o_1
XU$$1296 U$$1296/A U$$1328/B VGND VGND VPWR VPWR U$$1296/X sky130_fd_sc_hd__xor2_1
XFILLER_148_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_91_0 dadda_fa_5_91_0/A dadda_fa_5_91_0/B dadda_fa_5_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_92_0/A dadda_fa_6_91_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1090 final_adder.U$$188/A final_adder.U$$897/X VGND VGND VPWR VPWR
+ output347/A sky130_fd_sc_hd__xor2_1
XFILLER_144_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout804 U$$2667/B2 VGND VGND VPWR VPWR U$$2665/B2 sky130_fd_sc_hd__buf_4
Xfanout815 fanout820/X VGND VGND VPWR VPWR U$$2578/B2 sky130_fd_sc_hd__buf_2
Xdadda_fa_1_76_6 U$$3883/X U$$4016/X U$$4149/X VGND VGND VPWR VPWR dadda_fa_2_77_2/B
+ dadda_fa_2_76_5/B sky130_fd_sc_hd__fa_1
Xfanout826 U$$2463/B2 VGND VGND VPWR VPWR U$$2413/B2 sky130_fd_sc_hd__buf_4
Xfanout837 U$$2139/B2 VGND VGND VPWR VPWR U$$2097/B2 sky130_fd_sc_hd__buf_4
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout848 U$$2022/B2 VGND VGND VPWR VPWR U$$2014/B2 sky130_fd_sc_hd__buf_4
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout859 U$$1915/B2 VGND VGND VPWR VPWR U$$1911/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_140_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_5 U$$4401/X input222/X dadda_fa_1_69_5/CIN VGND VGND VPWR VPWR dadda_fa_2_70_2/A
+ dadda_fa_2_69_5/A sky130_fd_sc_hd__fa_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_96_0 dadda_ha_1_96_0/A U$$2327/X VGND VGND VPWR VPWR dadda_fa_3_97_0/A
+ dadda_fa_3_96_0/A sky130_fd_sc_hd__ha_1
XFILLER_6_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_100_1 dadda_fa_3_100_1/A dadda_fa_3_100_1/B dadda_fa_3_100_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_101_0/CIN dadda_fa_4_100_2/A sky130_fd_sc_hd__fa_1
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_121_0 dadda_fa_6_121_0/A dadda_fa_6_121_0/B dadda_fa_6_121_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_122_0/B dadda_fa_7_121_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_64_4 U$$1731/X U$$1864/X U$$1997/X VGND VGND VPWR VPWR dadda_fa_1_65_6/CIN
+ dadda_fa_1_64_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_41_3 dadda_fa_3_41_3/A dadda_fa_3_41_3/B dadda_fa_3_41_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_1/B dadda_fa_4_41_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$460 final_adder.U$$464/B final_adder.U$$460/B VGND VGND VPWR VPWR
+ final_adder.U$$584/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$471 final_adder.U$$470/B final_adder.U$$349/X final_adder.U$$345/X
+ VGND VGND VPWR VPWR final_adder.U$$471/X sky130_fd_sc_hd__a21o_1
XFILLER_17_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$310 U$$447/A1 U$$340/A2 U$$447/B1 U$$340/B2 VGND VGND VPWR VPWR U$$311/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$482 final_adder.U$$486/B final_adder.U$$482/B VGND VGND VPWR VPWR
+ final_adder.U$$606/B sky130_fd_sc_hd__and2_1
XU$$321 U$$321/A U$$353/B VGND VGND VPWR VPWR U$$321/X sky130_fd_sc_hd__xor2_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_34_2 dadda_fa_3_34_2/A dadda_fa_3_34_2/B dadda_fa_3_34_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_1/A dadda_fa_4_34_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$493 final_adder.U$$492/B final_adder.U$$371/X final_adder.U$$367/X
+ VGND VGND VPWR VPWR final_adder.U$$493/X sky130_fd_sc_hd__a21o_1
XU$$332 U$$58/A1 U$$362/A2 U$$60/A1 U$$362/B2 VGND VGND VPWR VPWR U$$333/A sky130_fd_sc_hd__a22o_1
XFILLER_17_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$343 U$$343/A U$$347/B VGND VGND VPWR VPWR U$$343/X sky130_fd_sc_hd__xor2_1
XU$$354 U$$902/A1 U$$362/A2 U$$902/B1 U$$362/B2 VGND VGND VPWR VPWR U$$355/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_27_1 U$$1524/X U$$1657/X U$$1790/X VGND VGND VPWR VPWR dadda_fa_4_28_0/CIN
+ dadda_fa_4_27_2/A sky130_fd_sc_hd__fa_1
XFILLER_17_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$365 U$$365/A U$$407/B VGND VGND VPWR VPWR U$$365/X sky130_fd_sc_hd__xor2_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$376 U$$650/A1 U$$386/A2 U$$650/B1 U$$386/B2 VGND VGND VPWR VPWR U$$377/A sky130_fd_sc_hd__a22o_1
XU$$387 U$$387/A U$$387/B VGND VGND VPWR VPWR U$$387/X sky130_fd_sc_hd__xor2_1
XU$$398 U$$672/A1 U$$406/A2 U$$672/B1 U$$406/B2 VGND VGND VPWR VPWR U$$399/A sky130_fd_sc_hd__a22o_1
XFILLER_158_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_86_5 dadda_fa_2_86_5/A dadda_fa_2_86_5/B dadda_fa_2_86_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_87_2/A dadda_fa_4_86_0/A sky130_fd_sc_hd__fa_2
XFILLER_114_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_79_4 dadda_fa_2_79_4/A dadda_fa_2_79_4/B dadda_fa_2_79_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_1/CIN dadda_fa_3_79_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1060 U$$1060/A U$$1062/B VGND VGND VPWR VPWR U$$1060/X sky130_fd_sc_hd__xor2_1
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1071 U$$934/A1 U$$1075/A2 U$$936/A1 U$$1075/B2 VGND VGND VPWR VPWR U$$1072/A sky130_fd_sc_hd__a22o_1
XU$$1082 U$$1082/A U$$1088/B VGND VGND VPWR VPWR U$$1082/X sky130_fd_sc_hd__xor2_1
XFILLER_148_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1093 U$$956/A1 U$$1093/A2 U$$1093/B1 U$$1093/B2 VGND VGND VPWR VPWR U$$1094/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_116_1 dadda_fa_5_116_1/A dadda_fa_5_116_1/B dadda_fa_5_116_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_117_0/B dadda_fa_7_116_0/A sky130_fd_sc_hd__fa_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_109_0 dadda_fa_5_109_0/A dadda_fa_5_109_0/B dadda_fa_5_109_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_110_0/A dadda_fa_6_109_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_81_4 U$$2829/X U$$2962/X U$$3095/X VGND VGND VPWR VPWR dadda_fa_2_82_2/B
+ dadda_fa_2_81_5/A sky130_fd_sc_hd__fa_1
XFILLER_132_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout601 U$$1891/A2 VGND VGND VPWR VPWR U$$1915/A2 sky130_fd_sc_hd__buf_6
XFILLER_137_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout612 U$$1593/A2 VGND VGND VPWR VPWR U$$1563/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout623 U$$259/A2 VGND VGND VPWR VPWR U$$271/A2 sky130_fd_sc_hd__buf_4
XFILLER_132_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_74_3 U$$2948/X U$$3081/X U$$3214/X VGND VGND VPWR VPWR dadda_fa_2_75_1/B
+ dadda_fa_2_74_4/B sky130_fd_sc_hd__fa_1
Xfanout634 U$$1502/A2 VGND VGND VPWR VPWR U$$1504/A2 sky130_fd_sc_hd__buf_6
Xfanout645 U$$1194/A2 VGND VGND VPWR VPWR U$$1164/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_51_2 dadda_fa_4_51_2/A dadda_fa_4_51_2/B dadda_fa_4_51_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_52_0/CIN dadda_fa_5_51_1/CIN sky130_fd_sc_hd__fa_1
Xfanout656 U$$981/B2 VGND VGND VPWR VPWR U$$979/B2 sky130_fd_sc_hd__buf_4
Xfanout667 U$$827/X VGND VGND VPWR VPWR U$$952/B2 sky130_fd_sc_hd__buf_8
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_2 U$$3333/X U$$3466/X U$$3599/X VGND VGND VPWR VPWR dadda_fa_2_68_1/A
+ dadda_fa_2_67_4/A sky130_fd_sc_hd__fa_1
XFILLER_85_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout678 U$$676/B2 VGND VGND VPWR VPWR U$$674/B2 sky130_fd_sc_hd__buf_4
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout689 U$$4369/B2 VGND VGND VPWR VPWR U$$4359/B2 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_4_44_1 dadda_fa_4_44_1/A dadda_fa_4_44_1/B dadda_fa_4_44_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_45_0/B dadda_fa_5_44_1/B sky130_fd_sc_hd__fa_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1002 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_21_0 dadda_fa_7_21_0/A dadda_fa_7_21_0/B dadda_fa_7_21_0/CIN VGND VGND
+ VPWR VPWR _318_/D _189_/D sky130_fd_sc_hd__fa_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_37_0 dadda_fa_4_37_0/A dadda_fa_4_37_0/B dadda_fa_4_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_38_0/A dadda_fa_5_37_1/A sky130_fd_sc_hd__fa_1
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_340_ _344_/CLK _340_/D VGND VGND VPWR VPWR _340_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_271_ _402_/CLK _271_/D VGND VGND VPWR VPWR _271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_70_4 U$$2009/X U$$2142/X VGND VGND VPWR VPWR dadda_fa_1_71_7/CIN dadda_fa_2_70_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_89_3 dadda_fa_3_89_3/A dadda_fa_3_89_3/B dadda_fa_3_89_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_1/B dadda_fa_4_89_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_56_2 U$$917/X U$$1050/X VGND VGND VPWR VPWR dadda_fa_1_57_8/A dadda_fa_2_56_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_111_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$6_1910 VGND VGND VPWR VPWR U$$6_1910/HI U$$6/A1 sky130_fd_sc_hd__conb_1
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_62_1 U$$530/X U$$663/X U$$796/X VGND VGND VPWR VPWR dadda_fa_1_63_5/CIN
+ dadda_fa_1_62_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3902 U$$4176/A1 U$$3906/A2 U$$4176/B1 U$$3906/B2 VGND VGND VPWR VPWR U$$3903/A
+ sky130_fd_sc_hd__a22o_1
XU$$4388_1840 VGND VGND VPWR VPWR U$$4388_1840/HI U$$4388/A2 sky130_fd_sc_hd__conb_1
XFILLER_134_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3913 U$$3913/A U$$3973/A VGND VGND VPWR VPWR U$$3913/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_55_0 U$$117/X U$$250/X U$$383/X VGND VGND VPWR VPWR dadda_fa_1_56_7/CIN
+ dadda_fa_1_55_8/CIN sky130_fd_sc_hd__fa_1
XU$$3924 U$$4196/B1 U$$3924/A2 U$$4198/B1 U$$3924/B2 VGND VGND VPWR VPWR U$$3925/A
+ sky130_fd_sc_hd__a22o_1
XU$$3935 U$$3935/A U$$3961/B VGND VGND VPWR VPWR U$$3935/X sky130_fd_sc_hd__xor2_1
XFILLER_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3946 U$$4081/B1 U$$3948/A2 U$$3948/A1 U$$3948/B2 VGND VGND VPWR VPWR U$$3947/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3957 U$$3957/A U$$3965/B VGND VGND VPWR VPWR U$$3957/X sky130_fd_sc_hd__xor2_1
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$290 final_adder.U$$292/B final_adder.U$$290/B VGND VGND VPWR VPWR
+ final_adder.U$$416/B sky130_fd_sc_hd__and2_1
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$140 U$$274/A U$$140/B VGND VGND VPWR VPWR U$$140/X sky130_fd_sc_hd__and2_1
XU$$3968 U$$4240/B1 U$$3970/A2 U$$4107/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3969/A
+ sky130_fd_sc_hd__a22o_1
XU$$3979 U$$3979/A1 U$$4005/A2 U$$3979/B1 U$$4005/B2 VGND VGND VPWR VPWR U$$3980/A
+ sky130_fd_sc_hd__a22o_1
XU$$151 U$$14/A1 U$$179/A2 U$$16/A1 U$$179/B2 VGND VGND VPWR VPWR U$$152/A sky130_fd_sc_hd__a22o_1
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$162 U$$162/A U$$214/B VGND VGND VPWR VPWR U$$162/X sky130_fd_sc_hd__xor2_1
XU$$173 U$$36/A1 U$$207/A2 U$$38/A1 U$$207/B2 VGND VGND VPWR VPWR U$$174/A sky130_fd_sc_hd__a22o_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$184 U$$184/A U$$220/B VGND VGND VPWR VPWR U$$184/X sky130_fd_sc_hd__xor2_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$195 U$$58/A1 U$$229/A2 U$$60/A1 U$$229/B2 VGND VGND VPWR VPWR U$$196/A sky130_fd_sc_hd__a22o_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_91_3 U$$4312/X U$$4445/X input247/X VGND VGND VPWR VPWR dadda_fa_3_92_1/B
+ dadda_fa_3_91_3/B sky130_fd_sc_hd__fa_1
XFILLER_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_84_2 dadda_fa_2_84_2/A dadda_fa_2_84_2/B dadda_fa_2_84_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_1/A dadda_fa_3_84_3/A sky130_fd_sc_hd__fa_1
Xoutput259 output259/A VGND VGND VPWR VPWR o[101] sky130_fd_sc_hd__buf_2
XFILLER_88_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_61_1 dadda_fa_5_61_1/A dadda_fa_5_61_1/B dadda_fa_5_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_62_0/B dadda_fa_7_61_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_77_1 dadda_fa_2_77_1/A dadda_fa_2_77_1/B dadda_fa_2_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_0/CIN dadda_fa_3_77_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_54_0 dadda_fa_5_54_0/A dadda_fa_5_54_0/B dadda_fa_5_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_55_0/A dadda_fa_6_54_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_53_8 U$$3571/X input205/X dadda_fa_1_53_8/CIN VGND VGND VPWR VPWR dadda_fa_2_54_3/A
+ dadda_fa_3_53_0/A sky130_fd_sc_hd__fa_1
XFILLER_49_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_100_0 dadda_fa_2_100_0/A U$$2601/X U$$2734/X VGND VGND VPWR VPWR dadda_fa_3_101_1/B
+ dadda_fa_3_100_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_24_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_99_2 dadda_fa_4_99_2/A dadda_fa_4_99_2/B dadda_fa_4_99_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_100_0/CIN dadda_fa_5_99_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1239_1784 VGND VGND VPWR VPWR U$$1239_1784/HI U$$1239/A1 sky130_fd_sc_hd__conb_1
Xdadda_fa_7_69_0 dadda_fa_7_69_0/A dadda_fa_7_69_0/B dadda_fa_7_69_0/CIN VGND VGND
+ VPWR VPWR _366_/D _237_/D sky130_fd_sc_hd__fa_1
XFILLER_155_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1407 U$$2745/A2 VGND VGND VPWR VPWR U$$2724/B sky130_fd_sc_hd__buf_4
Xfanout1418 fanout1419/X VGND VGND VPWR VPWR U$$2602/A sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_1_72_0 U$$2013/X U$$2146/X U$$2279/X VGND VGND VPWR VPWR dadda_fa_2_73_0/B
+ dadda_fa_2_72_3/B sky130_fd_sc_hd__fa_1
Xfanout420 U$$4369/A2 VGND VGND VPWR VPWR U$$4349/A2 sky130_fd_sc_hd__buf_4
Xfanout431 U$$545/A2 VGND VGND VPWR VPWR U$$505/A2 sky130_fd_sc_hd__buf_4
XFILLER_24_1003 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1429 U$$2402/B VGND VGND VPWR VPWR U$$2396/B sky130_fd_sc_hd__buf_6
Xfanout442 U$$102/A2 VGND VGND VPWR VPWR U$$86/A2 sky130_fd_sc_hd__buf_4
Xfanout453 U$$3977/X VGND VGND VPWR VPWR U$$4043/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1011 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout464 U$$3966/A2 VGND VGND VPWR VPWR U$$3948/A2 sky130_fd_sc_hd__buf_4
XFILLER_48_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout475 U$$3703/X VGND VGND VPWR VPWR U$$3833/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout486 U$$3473/A2 VGND VGND VPWR VPWR U$$3511/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout497 U$$3306/A2 VGND VGND VPWR VPWR U$$3390/A2 sky130_fd_sc_hd__buf_6
XU$$3209 U$$878/B1 U$$3255/A2 U$$745/A1 U$$3255/B2 VGND VGND VPWR VPWR U$$3210/A sky130_fd_sc_hd__a22o_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2508 U$$2780/B1 U$$2548/A2 U$$2647/A1 U$$2548/B2 VGND VGND VPWR VPWR U$$2509/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2519 U$$2519/A U$$2541/B VGND VGND VPWR VPWR U$$2519/X sky130_fd_sc_hd__xor2_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1807 U$$26/A1 U$$1881/A2 U$$28/A1 U$$1881/B2 VGND VGND VPWR VPWR U$$1808/A sky130_fd_sc_hd__a22o_1
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1818 U$$1818/A U$$1832/B VGND VGND VPWR VPWR U$$1818/X sky130_fd_sc_hd__xor2_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1829 U$$596/A1 U$$1829/A2 U$$596/B1 U$$1829/B2 VGND VGND VPWR VPWR U$$1830/A sky130_fd_sc_hd__a22o_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_323_ _328_/CLK _323_/D VGND VGND VPWR VPWR _323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_254_ _382_/CLK _254_/D VGND VGND VPWR VPWR _254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_185_ _321_/CLK _185_/D VGND VGND VPWR VPWR _185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_94_1 dadda_fa_3_94_1/A dadda_fa_3_94_1/B dadda_fa_3_94_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_0/CIN dadda_fa_4_94_2/A sky130_fd_sc_hd__fa_1
XFILLER_171_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_71_0 dadda_fa_6_71_0/A dadda_fa_6_71_0/B dadda_fa_6_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_72_0/B dadda_fa_7_71_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_87_0 dadda_fa_3_87_0/A dadda_fa_3_87_0/B dadda_fa_3_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_0/B dadda_fa_4_87_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_123_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4400 U$$4400/A1 U$$4388/X U$$4400/B1 U$$4428/B2 VGND VGND VPWR VPWR U$$4401/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4411 U$$4411/A U$$4411/B VGND VGND VPWR VPWR U$$4411/X sky130_fd_sc_hd__xor2_1
XU$$4422 U$$4422/A1 U$$4388/X U$$4424/A1 U$$4508/B2 VGND VGND VPWR VPWR U$$4423/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4433 U$$4433/A U$$4433/B VGND VGND VPWR VPWR U$$4433/X sky130_fd_sc_hd__xor2_1
XFILLER_64_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4444 U$$4444/A1 U$$4388/X U$$4446/A1 U$$4506/B2 VGND VGND VPWR VPWR U$$4445/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4455 U$$4455/A U$$4455/B VGND VGND VPWR VPWR U$$4455/X sky130_fd_sc_hd__xor2_1
XU$$3710 U$$3710/A U$$3790/B VGND VGND VPWR VPWR U$$3710/X sky130_fd_sc_hd__xor2_1
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3721 U$$4132/A1 U$$3757/A2 U$$4132/B1 U$$3757/B2 VGND VGND VPWR VPWR U$$3722/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_49_5 dadda_fa_2_49_5/A dadda_fa_2_49_5/B dadda_fa_2_49_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_2/A dadda_fa_4_49_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_4_116_0 U$$3830/X U$$3963/X U$$4096/X VGND VGND VPWR VPWR dadda_fa_5_117_0/A
+ dadda_fa_5_116_1/A sky130_fd_sc_hd__fa_1
XU$$4466 U$$4466/A1 U$$4388/X U$$4468/A1 U$$4488/B2 VGND VGND VPWR VPWR U$$4467/A
+ sky130_fd_sc_hd__a22o_1
XU$$3732 U$$3732/A U$$3734/B VGND VGND VPWR VPWR U$$3732/X sky130_fd_sc_hd__xor2_1
XU$$4477 U$$4477/A U$$4477/B VGND VGND VPWR VPWR U$$4477/X sky130_fd_sc_hd__xor2_1
XFILLER_65_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4488 U$$4488/A1 U$$4388/X U$$4490/A1 U$$4488/B2 VGND VGND VPWR VPWR U$$4489/A
+ sky130_fd_sc_hd__a22o_1
XU$$3743 U$$4152/B1 U$$3791/A2 U$$4017/B1 U$$3791/B2 VGND VGND VPWR VPWR U$$3744/A
+ sky130_fd_sc_hd__a22o_1
XU$$3754 U$$3754/A U$$3836/A VGND VGND VPWR VPWR U$$3754/X sky130_fd_sc_hd__xor2_1
XU$$4499 U$$4499/A U$$4499/B VGND VGND VPWR VPWR U$$4499/X sky130_fd_sc_hd__xor2_1
XU$$3765 U$$4176/A1 U$$3773/A2 U$$4176/B1 U$$3773/B2 VGND VGND VPWR VPWR U$$3766/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3776 U$$3776/A U$$3836/A VGND VGND VPWR VPWR U$$3776/X sky130_fd_sc_hd__xor2_1
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3787 U$$910/A1 U$$3791/A2 U$$912/A1 U$$3791/B2 VGND VGND VPWR VPWR U$$3788/A sky130_fd_sc_hd__a22o_1
XU$$3798 U$$3798/A U$$3816/B VGND VGND VPWR VPWR U$$3798/X sky130_fd_sc_hd__xor2_1
XFILLER_33_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1778_1793 VGND VGND VPWR VPWR U$$1778_1793/HI U$$1778/B1 sky130_fd_sc_hd__conb_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_51_5 U$$2104/X U$$2237/X U$$2370/X VGND VGND VPWR VPWR dadda_fa_2_52_2/A
+ dadda_fa_2_51_5/A sky130_fd_sc_hd__fa_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$909 U$$909/A U$$913/B VGND VGND VPWR VPWR U$$909/X sky130_fd_sc_hd__xor2_1
XFILLER_141_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_44_4 U$$1691/X U$$1824/X U$$1957/X VGND VGND VPWR VPWR dadda_fa_2_45_3/CIN
+ dadda_fa_2_44_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_14_2 U$$980/B input162/X dadda_ha_3_14_0/SUM VGND VGND VPWR VPWR dadda_fa_5_15_0/CIN
+ dadda_fa_5_14_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_93_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1204 U$$3870/A1 VGND VGND VPWR VPWR U$$854/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout1215 U$$3181/B1 VGND VGND VPWR VPWR U$$32/A1 sky130_fd_sc_hd__buf_4
Xfanout1226 U$$2631/A1 VGND VGND VPWR VPWR U$$850/A1 sky130_fd_sc_hd__buf_4
Xfanout1237 input65/X VGND VGND VPWR VPWR U$$3981/A1 sky130_fd_sc_hd__buf_4
XFILLER_94_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1248 U$$639/B VGND VGND VPWR VPWR U$$643/B sky130_fd_sc_hd__clkbuf_4
Xfanout1259 U$$547/A VGND VGND VPWR VPWR U$$522/B sky130_fd_sc_hd__buf_8
XFILLER_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3006 U$$3006/A U$$3013/A VGND VGND VPWR VPWR U$$3006/X sky130_fd_sc_hd__xor2_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3017 U$$3151/A U$$3017/B VGND VGND VPWR VPWR U$$3017/X sky130_fd_sc_hd__and2_1
XFILLER_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3028 U$$3163/B1 U$$3066/A2 U$$3030/A1 U$$3066/B2 VGND VGND VPWR VPWR U$$3029/A
+ sky130_fd_sc_hd__a22o_1
XU$$3039 U$$3039/A U$$3077/B VGND VGND VPWR VPWR U$$3039/X sky130_fd_sc_hd__xor2_1
XU$$2305 U$$2305/A U$$2329/A VGND VGND VPWR VPWR U$$2305/X sky130_fd_sc_hd__xor2_1
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2316 U$$4234/A1 U$$2320/A2 U$$4234/B1 U$$2320/B2 VGND VGND VPWR VPWR U$$2317/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2327 U$$2327/A U$$2327/B VGND VGND VPWR VPWR U$$2327/X sky130_fd_sc_hd__xor2_1
XU$$2338 U$$2338/A U$$2412/B VGND VGND VPWR VPWR U$$2338/X sky130_fd_sc_hd__xor2_1
XFILLER_43_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1604 U$$1604/A U$$1608/B VGND VGND VPWR VPWR U$$1604/X sky130_fd_sc_hd__xor2_1
XU$$2349 U$$4404/A1 U$$2407/A2 U$$981/A1 U$$2407/B2 VGND VGND VPWR VPWR U$$2350/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1615 U$$654/B1 U$$1625/A2 U$$521/A1 U$$1625/B2 VGND VGND VPWR VPWR U$$1616/A sky130_fd_sc_hd__a22o_1
XFILLER_43_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1626 U$$1626/A U$$1626/B VGND VGND VPWR VPWR U$$1626/X sky130_fd_sc_hd__xor2_1
XFILLER_15_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1637 U$$4512/B1 U$$1641/A2 U$$4377/B1 U$$1641/B2 VGND VGND VPWR VPWR U$$1638/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1648 U$$1646/Y input17/X U$$1630/B U$$1647/X U$$1644/Y VGND VGND VPWR VPWR U$$1648/X
+ sky130_fd_sc_hd__a32o_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1659 U$$1659/A U$$1697/B VGND VGND VPWR VPWR U$$1659/X sky130_fd_sc_hd__xor2_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_306_ _319_/CLK _306_/D VGND VGND VPWR VPWR _306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_237_ _366_/CLK _237_/D VGND VGND VPWR VPWR _237_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_168_ _319_/CLK _168_/D VGND VGND VPWR VPWR _168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_61_4 dadda_fa_2_61_4/A dadda_fa_2_61_4/B dadda_fa_2_61_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_1/CIN dadda_fa_3_61_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1760 U$$914/B1 VGND VGND VPWR VPWR U$$3382/A1 sky130_fd_sc_hd__buf_6
Xfanout1771 U$$3376/B1 VGND VGND VPWR VPWR U$$90/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_54_3 dadda_fa_2_54_3/A dadda_fa_2_54_3/B dadda_fa_2_54_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_1/B dadda_fa_3_54_3/B sky130_fd_sc_hd__fa_1
XU$$4230 U$$4365/B1 U$$4236/A2 U$$4367/B1 U$$4236/B2 VGND VGND VPWR VPWR U$$4231/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4241 U$$4241/A U$$4241/B VGND VGND VPWR VPWR U$$4241/X sky130_fd_sc_hd__xor2_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4252 U$$4250/B U$$4247/A input59/X U$$4247/Y VGND VGND VPWR VPWR U$$4252/X sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_47_2 dadda_fa_2_47_2/A dadda_fa_2_47_2/B dadda_fa_2_47_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_1/A dadda_fa_3_47_3/A sky130_fd_sc_hd__fa_1
XU$$4263 U$$4400/A1 U$$4295/A2 U$$4400/B1 U$$4295/B2 VGND VGND VPWR VPWR U$$4264/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4274 U$$4274/A U$$4322/B VGND VGND VPWR VPWR U$$4274/X sky130_fd_sc_hd__xor2_1
XFILLER_66_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4285 U$$4420/B1 U$$4309/A2 U$$4287/A1 U$$4309/B2 VGND VGND VPWR VPWR U$$4286/A
+ sky130_fd_sc_hd__a22o_1
XU$$3540 U$$3540/A U$$3561/A VGND VGND VPWR VPWR U$$3540/X sky130_fd_sc_hd__xor2_1
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_24_1 dadda_fa_5_24_1/A dadda_fa_5_24_1/B dadda_fa_5_24_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_25_0/B dadda_fa_7_24_0/A sky130_fd_sc_hd__fa_2
XFILLER_80_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3551 U$$3551/A1 U$$3557/A2 U$$3964/A1 U$$3557/B2 VGND VGND VPWR VPWR U$$3552/A
+ sky130_fd_sc_hd__a22o_1
XU$$4296 U$$4296/A U$$4384/A VGND VGND VPWR VPWR U$$4296/X sky130_fd_sc_hd__xor2_1
XFILLER_37_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3562 U$$3562/A VGND VGND VPWR VPWR U$$3562/Y sky130_fd_sc_hd__inv_1
XU$$3573 U$$3573/A U$$3615/B VGND VGND VPWR VPWR U$$3573/X sky130_fd_sc_hd__xor2_1
XU$$3584 U$$4132/A1 U$$3604/A2 U$$4132/B1 U$$3604/B2 VGND VGND VPWR VPWR U$$3585/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_17_0 dadda_fa_5_17_0/A dadda_fa_5_17_0/B dadda_fa_5_17_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_18_0/A dadda_fa_6_17_0/CIN sky130_fd_sc_hd__fa_1
XU$$3595 U$$3595/A U$$3601/B VGND VGND VPWR VPWR U$$3595/X sky130_fd_sc_hd__xor2_1
XU$$2850 U$$4220/A1 U$$2874/A2 U$$4220/B1 U$$2874/B2 VGND VGND VPWR VPWR U$$2851/A
+ sky130_fd_sc_hd__a22o_1
XU$$2861 U$$2861/A U$$2871/B VGND VGND VPWR VPWR U$$2861/X sky130_fd_sc_hd__xor2_1
XFILLER_34_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2872 U$$3692/B1 U$$2872/A2 U$$3559/A1 U$$2872/B2 VGND VGND VPWR VPWR U$$2873/A
+ sky130_fd_sc_hd__a22o_1
XU$$2883 U$$2883/A1 U$$2929/A2 U$$3022/A1 U$$2929/B2 VGND VGND VPWR VPWR U$$2884/A
+ sky130_fd_sc_hd__a22o_1
XU$$2894 U$$2894/A U$$2926/B VGND VGND VPWR VPWR U$$2894/X sky130_fd_sc_hd__xor2_1
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$801 final_adder.U$$800/B final_adder.U$$721/X final_adder.U$$689/X
+ VGND VGND VPWR VPWR final_adder.U$$801/X sky130_fd_sc_hd__a21o_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$823 final_adder.U$$790/A final_adder.U$$623/X final_adder.U$$711/X
+ VGND VGND VPWR VPWR final_adder.U$$823/X sky130_fd_sc_hd__a21o_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$845 final_adder.U$$748/X final_adder.U$$813/X final_adder.U$$749/X
+ VGND VGND VPWR VPWR final_adder.U$$845/X sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$867 final_adder.U$$770/X final_adder.U$$723/X final_adder.U$$771/X
+ VGND VGND VPWR VPWR final_adder.U$$867/X sky130_fd_sc_hd__a21o_1
XU$$706 U$$706/A U$$774/B VGND VGND VPWR VPWR U$$706/X sky130_fd_sc_hd__xor2_1
XU$$717 U$$991/A1 U$$763/A2 U$$993/A1 U$$763/B2 VGND VGND VPWR VPWR U$$718/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$889 final_adder.U$$792/X final_adder.U$$625/X final_adder.U$$793/X
+ VGND VGND VPWR VPWR final_adder.U$$889/X sky130_fd_sc_hd__a21o_1
XU$$728 U$$728/A U$$764/B VGND VGND VPWR VPWR U$$728/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_42_1 U$$490/X U$$623/X U$$756/X VGND VGND VPWR VPWR dadda_fa_2_43_3/B
+ dadda_fa_2_42_5/A sky130_fd_sc_hd__fa_1
XFILLER_44_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$739 U$$739/A1 U$$819/A2 U$$741/A1 U$$819/B2 VGND VGND VPWR VPWR U$$740/A sky130_fd_sc_hd__a22o_1
XFILLER_45_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_71_3 dadda_fa_3_71_3/A dadda_fa_3_71_3/B dadda_fa_3_71_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_1/B dadda_fa_4_71_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1001 fanout999/A VGND VGND VPWR VPWR U$$4460/A1 sky130_fd_sc_hd__buf_2
Xfanout1012 U$$70/B1 VGND VGND VPWR VPWR U$$894/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_64_2 dadda_fa_3_64_2/A dadda_fa_3_64_2/B dadda_fa_3_64_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_1/A dadda_fa_4_64_2/B sky130_fd_sc_hd__fa_1
Xfanout1023 U$$1189/B VGND VGND VPWR VPWR U$$1231/B sky130_fd_sc_hd__clkbuf_4
Xfanout1034 U$$4315/B1 VGND VGND VPWR VPWR U$$4043/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1045 U$$4257/B1 VGND VGND VPWR VPWR U$$2887/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1056 U$$612/B1 VGND VGND VPWR VPWR U$$749/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_57_1 dadda_fa_3_57_1/A dadda_fa_3_57_1/B dadda_fa_3_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_0/CIN dadda_fa_4_57_2/A sky130_fd_sc_hd__fa_1
XFILLER_120_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1067 U$$4446/B1 VGND VGND VPWR VPWR U$$3763/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout1078 U$$469/B1 VGND VGND VPWR VPWR U$$60/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_34_0 dadda_fa_6_34_0/A dadda_fa_6_34_0/B dadda_fa_6_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_35_0/B dadda_fa_7_34_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1089 U$$878/B1 VGND VGND VPWR VPWR U$$880/A1 sky130_fd_sc_hd__buf_4
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2102 U$$2102/A U$$2106/B VGND VGND VPWR VPWR U$$2102/X sky130_fd_sc_hd__xor2_1
XU$$2113 U$$880/A1 U$$2147/A2 U$$882/A1 U$$2147/B2 VGND VGND VPWR VPWR U$$2114/A sky130_fd_sc_hd__a22o_1
XU$$2124 U$$2124/A U$$2130/B VGND VGND VPWR VPWR U$$2124/X sky130_fd_sc_hd__xor2_1
XU$$2135 U$$902/A1 U$$2139/A2 U$$902/B1 U$$2139/B2 VGND VGND VPWR VPWR U$$2136/A sky130_fd_sc_hd__a22o_1
XFILLER_63_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1401 U$$1401/A U$$1415/B VGND VGND VPWR VPWR U$$1401/X sky130_fd_sc_hd__xor2_1
XU$$2146 U$$2146/A U$$2148/B VGND VGND VPWR VPWR U$$2146/X sky130_fd_sc_hd__xor2_1
XFILLER_62_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2157 U$$4486/A1 U$$2181/A2 U$$4486/B1 U$$2181/B2 VGND VGND VPWR VPWR U$$2158/A
+ sky130_fd_sc_hd__a22o_1
XU$$1412 U$$40/B1 U$$1414/A2 U$$316/B1 U$$1414/B2 VGND VGND VPWR VPWR U$$1413/A sky130_fd_sc_hd__a22o_1
XFILLER_34_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1423 U$$1423/A U$$1427/B VGND VGND VPWR VPWR U$$1423/X sky130_fd_sc_hd__xor2_1
XU$$2168 U$$2168/A U$$2168/B VGND VGND VPWR VPWR U$$2168/X sky130_fd_sc_hd__xor2_1
XU$$1434 U$$884/B1 U$$1460/A2 U$$64/B1 U$$1460/B2 VGND VGND VPWR VPWR U$$1435/A sky130_fd_sc_hd__a22o_1
XU$$2179 U$$2862/B1 U$$2189/A2 U$$2179/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2180/A
+ sky130_fd_sc_hd__a22o_1
XU$$1445 U$$1445/A U$$1449/B VGND VGND VPWR VPWR U$$1445/X sky130_fd_sc_hd__xor2_1
XU$$1456 U$$632/B1 U$$1460/A2 U$$499/A1 U$$1460/B2 VGND VGND VPWR VPWR U$$1457/A sky130_fd_sc_hd__a22o_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1467 U$$1467/A U$$1507/A VGND VGND VPWR VPWR U$$1467/X sky130_fd_sc_hd__xor2_1
XU$$1478 U$$654/B1 U$$1480/A2 U$$521/A1 U$$1480/B2 VGND VGND VPWR VPWR U$$1479/A sky130_fd_sc_hd__a22o_1
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1489 U$$1489/A U$$1491/B VGND VGND VPWR VPWR U$$1489/X sky130_fd_sc_hd__xor2_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_866 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_107_0 dadda_fa_7_107_0/A dadda_fa_7_107_0/B dadda_fa_7_107_0/CIN VGND
+ VGND VPWR VPWR _404_/D _275_/D sky130_fd_sc_hd__fa_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_941 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$108 _404_/Q _276_/Q VGND VGND VPWR VPWR final_adder.U$$917/B1 final_adder.U$$146/A
+ sky130_fd_sc_hd__ha_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$119 _415_/Q _287_/Q VGND VGND VPWR VPWR final_adder.U$$137/B1 final_adder.U$$136/B
+ sky130_fd_sc_hd__ha_2
Xdadda_fa_2_52_0 dadda_fa_2_52_0/A dadda_fa_2_52_0/B dadda_fa_2_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_0/B dadda_fa_3_52_2/B sky130_fd_sc_hd__fa_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1590 U$$121/B VGND VGND VPWR VPWR U$$77/B sky130_fd_sc_hd__buf_6
XFILLER_39_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4060 U$$4060/A U$$4082/B VGND VGND VPWR VPWR U$$4060/X sky130_fd_sc_hd__xor2_1
XU$$4071 U$$4482/A1 U$$4093/A2 U$$4484/A1 U$$4093/B2 VGND VGND VPWR VPWR U$$4072/A
+ sky130_fd_sc_hd__a22o_1
XU$$4082 U$$4082/A U$$4082/B VGND VGND VPWR VPWR U$$4082/X sky130_fd_sc_hd__xor2_1
XU$$4093 U$$4093/A1 U$$4093/A2 U$$4093/B1 U$$4093/B2 VGND VGND VPWR VPWR U$$4094/A
+ sky130_fd_sc_hd__a22o_1
XU$$3370 U$$3370/A1 U$$3372/A2 U$$3370/B1 U$$3372/B2 VGND VGND VPWR VPWR U$$3371/A
+ sky130_fd_sc_hd__a22o_1
XU$$3381 U$$3381/A U$$3424/A VGND VGND VPWR VPWR U$$3381/X sky130_fd_sc_hd__xor2_1
XU$$3392 U$$4349/B1 U$$3416/A2 U$$4214/B1 U$$3416/B2 VGND VGND VPWR VPWR U$$3393/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2680 U$$2680/A U$$2724/B VGND VGND VPWR VPWR U$$2680/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_6_0 U$$19/X U$$152/X U$$285/X VGND VGND VPWR VPWR dadda_fa_6_7_0/A dadda_fa_6_6_0/CIN
+ sky130_fd_sc_hd__fa_1
XU$$2691 U$$3376/A1 U$$2711/A2 U$$3376/B1 U$$2711/B2 VGND VGND VPWR VPWR U$$2692/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1990 U$$70/B1 U$$2006/A2 U$$620/B1 U$$2006/B2 VGND VGND VPWR VPWR U$$1991/A sky130_fd_sc_hd__a22o_1
XFILLER_22_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_81_2 dadda_fa_4_81_2/A dadda_fa_4_81_2/B dadda_fa_4_81_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_82_0/CIN dadda_fa_5_81_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_4_118_0_1939 VGND VGND VPWR VPWR dadda_fa_4_118_0/A dadda_fa_4_118_0_1939/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_116_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_74_1 dadda_fa_4_74_1/A dadda_fa_4_74_1/B dadda_fa_4_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_75_0/B dadda_fa_5_74_1/B sky130_fd_sc_hd__fa_1
XFILLER_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_51_0 dadda_fa_7_51_0/A dadda_fa_7_51_0/B dadda_fa_7_51_0/CIN VGND VGND
+ VPWR VPWR _348_/D _219_/D sky130_fd_sc_hd__fa_1
XFILLER_103_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_67_0 dadda_fa_4_67_0/A dadda_fa_4_67_0/B dadda_fa_4_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_68_0/A dadda_fa_5_67_1/A sky130_fd_sc_hd__fa_1
XFILLER_0_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput104 b[45] VGND VGND VPWR VPWR input104/X sky130_fd_sc_hd__buf_4
Xinput115 b[55] VGND VGND VPWR VPWR input115/X sky130_fd_sc_hd__buf_2
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput126 b[7] VGND VGND VPWR VPWR input126/X sky130_fd_sc_hd__buf_2
Xinput137 c[107] VGND VGND VPWR VPWR input137/X sky130_fd_sc_hd__clkbuf_4
XFILLER_102_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput148 c[117] VGND VGND VPWR VPWR input148/X sky130_fd_sc_hd__buf_2
Xinput159 c[127] VGND VGND VPWR VPWR input159/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$631 final_adder.U$$630/B final_adder.U$$527/X final_adder.U$$511/X
+ VGND VGND VPWR VPWR final_adder.U$$631/X sky130_fd_sc_hd__a21o_1
XFILLER_5_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$642 final_adder.U$$658/B final_adder.U$$642/B VGND VGND VPWR VPWR
+ final_adder.U$$754/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$653 final_adder.U$$652/B final_adder.U$$549/X final_adder.U$$533/X
+ VGND VGND VPWR VPWR final_adder.U$$653/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$664 final_adder.U$$680/B final_adder.U$$664/B VGND VGND VPWR VPWR
+ final_adder.U$$776/B sky130_fd_sc_hd__and2_1
XU$$503 U$$503/A1 U$$543/A2 U$$505/A1 U$$543/B2 VGND VGND VPWR VPWR U$$504/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$675 final_adder.U$$674/B final_adder.U$$571/X final_adder.U$$555/X
+ VGND VGND VPWR VPWR final_adder.U$$675/X sky130_fd_sc_hd__a21o_1
XU$$514 U$$514/A U$$522/B VGND VGND VPWR VPWR U$$514/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$686 final_adder.U$$702/B final_adder.U$$686/B VGND VGND VPWR VPWR
+ final_adder.U$$798/B sky130_fd_sc_hd__and2_1
XFILLER_29_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$525 U$$936/A1 U$$539/A2 U$$936/B1 U$$539/B2 VGND VGND VPWR VPWR U$$526/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$697 final_adder.U$$696/B final_adder.U$$593/X final_adder.U$$577/X
+ VGND VGND VPWR VPWR final_adder.U$$697/X sky130_fd_sc_hd__a21o_1
XU$$536 U$$536/A U$$536/B VGND VGND VPWR VPWR U$$536/X sky130_fd_sc_hd__xor2_1
XU$$547 U$$547/A VGND VGND VPWR VPWR U$$547/Y sky130_fd_sc_hd__inv_1
XU$$558 U$$8/B1 U$$610/A2 U$$12/A1 U$$610/B2 VGND VGND VPWR VPWR U$$559/A sky130_fd_sc_hd__a22o_1
XU$$569 U$$569/A U$$639/B VGND VGND VPWR VPWR U$$569/X sky130_fd_sc_hd__xor2_1
XFILLER_60_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_980 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1220 U$$946/A1 U$$1226/A2 U$$948/A1 U$$1226/B2 VGND VGND VPWR VPWR U$$1221/A sky130_fd_sc_hd__a22o_1
XU$$1231 U$$1231/A U$$1231/B VGND VGND VPWR VPWR U$$1231/X sky130_fd_sc_hd__xor2_1
XFILLER_62_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1242 U$$1242/A U$$1282/B VGND VGND VPWR VPWR U$$1242/X sky130_fd_sc_hd__xor2_1
XU$$1253 U$$2897/A1 U$$1327/A2 U$$2897/B1 U$$1327/B2 VGND VGND VPWR VPWR U$$1254/A
+ sky130_fd_sc_hd__a22o_1
XU$$1264 U$$1264/A U$$1300/B VGND VGND VPWR VPWR U$$1264/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_42_clk _218_/CLK VGND VGND VPWR VPWR _364_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1275 U$$42/A1 U$$1309/A2 U$$44/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1276/A sky130_fd_sc_hd__a22o_1
XU$$1286 U$$1286/A U$$1300/B VGND VGND VPWR VPWR U$$1286/X sky130_fd_sc_hd__xor2_1
XU$$1297 U$$64/A1 U$$1327/A2 U$$64/B1 U$$1327/B2 VGND VGND VPWR VPWR U$$1298/A sky130_fd_sc_hd__a22o_1
XFILLER_30_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_91_1 dadda_fa_5_91_1/A dadda_fa_5_91_1/B dadda_fa_5_91_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_92_0/B dadda_fa_7_91_0/A sky130_fd_sc_hd__fa_1
XFILLER_157_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_84_0 dadda_fa_5_84_0/A dadda_fa_5_84_0/B dadda_fa_5_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_85_0/A dadda_fa_6_84_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1080 final_adder.U$$198/A final_adder.U$$811/X VGND VGND VPWR VPWR
+ output336/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1091 final_adder.U$$188/B final_adder.U$$959/X VGND VGND VPWR VPWR
+ output348/A sky130_fd_sc_hd__xor2_1
XFILLER_104_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout805 U$$2608/X VGND VGND VPWR VPWR U$$2667/B2 sky130_fd_sc_hd__buf_4
XFILLER_131_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout816 fanout820/X VGND VGND VPWR VPWR U$$2546/B2 sky130_fd_sc_hd__buf_6
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout827 U$$2463/B2 VGND VGND VPWR VPWR U$$2459/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_76_7 U$$4282/X U$$4415/X input230/X VGND VGND VPWR VPWR dadda_fa_2_77_2/CIN
+ dadda_fa_2_76_5/CIN sky130_fd_sc_hd__fa_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout838 U$$2060/X VGND VGND VPWR VPWR U$$2139/B2 sky130_fd_sc_hd__clkbuf_8
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout849 U$$2052/B2 VGND VGND VPWR VPWR U$$2046/B2 sky130_fd_sc_hd__buf_4
XFILLER_86_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_6 dadda_fa_1_69_6/A dadda_fa_1_69_6/B dadda_fa_1_69_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_70_2/B dadda_fa_2_69_5/B sky130_fd_sc_hd__fa_1
XFILLER_85_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_969 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_clk _388_/CLK VGND VGND VPWR VPWR _383_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_99_0 dadda_fa_7_99_0/A dadda_fa_7_99_0/B dadda_fa_7_99_0/CIN VGND VGND
+ VPWR VPWR _396_/D _267_/D sky130_fd_sc_hd__fa_1
XFILLER_21_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_100_2 dadda_fa_3_100_2/A dadda_fa_3_100_2/B dadda_fa_3_100_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_101_1/A dadda_fa_4_100_2/B sky130_fd_sc_hd__fa_1
XFILLER_163_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_64_5 U$$2130/X U$$2263/X U$$2396/X VGND VGND VPWR VPWR dadda_fa_1_65_7/A
+ dadda_fa_2_64_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_6_114_0 dadda_fa_6_114_0/A dadda_fa_6_114_0/B dadda_fa_6_114_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_115_0/B dadda_fa_7_114_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_18_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$450 final_adder.U$$454/B final_adder.U$$450/B VGND VGND VPWR VPWR
+ final_adder.U$$574/B sky130_fd_sc_hd__and2_1
XFILLER_91_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$300 U$$26/A1 U$$340/A2 U$$28/A1 U$$340/B2 VGND VGND VPWR VPWR U$$301/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$461 final_adder.U$$460/B final_adder.U$$339/X final_adder.U$$335/X
+ VGND VGND VPWR VPWR final_adder.U$$461/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$472 final_adder.U$$476/B final_adder.U$$472/B VGND VGND VPWR VPWR
+ final_adder.U$$596/B sky130_fd_sc_hd__and2_1
XFILLER_17_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$311 U$$311/A U$$341/B VGND VGND VPWR VPWR U$$311/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$483 final_adder.U$$482/B final_adder.U$$361/X final_adder.U$$357/X
+ VGND VGND VPWR VPWR final_adder.U$$483/X sky130_fd_sc_hd__a21o_1
XU$$322 U$$868/B1 U$$352/A2 U$$735/A1 U$$352/B2 VGND VGND VPWR VPWR U$$323/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_34_3 dadda_fa_3_34_3/A dadda_fa_3_34_3/B dadda_fa_3_34_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_1/B dadda_fa_4_34_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$494 final_adder.U$$498/B final_adder.U$$494/B VGND VGND VPWR VPWR
+ final_adder.U$$610/A sky130_fd_sc_hd__and2_1
XU$$333 U$$333/A U$$363/B VGND VGND VPWR VPWR U$$333/X sky130_fd_sc_hd__xor2_1
XU$$344 U$$479/B1 U$$346/A2 U$$72/A1 U$$346/B2 VGND VGND VPWR VPWR U$$345/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_27_2 input176/X dadda_fa_3_27_2/B dadda_fa_3_27_2/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_28_1/A dadda_fa_4_27_2/B sky130_fd_sc_hd__fa_1
XU$$355 U$$355/A U$$363/B VGND VGND VPWR VPWR U$$355/X sky130_fd_sc_hd__xor2_1
XFILLER_83_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$366 U$$92/A1 U$$406/A2 U$$94/A1 U$$406/B2 VGND VGND VPWR VPWR U$$367/A sky130_fd_sc_hd__a22o_1
XFILLER_17_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$377 U$$377/A U$$387/B VGND VGND VPWR VPWR U$$377/X sky130_fd_sc_hd__xor2_1
XFILLER_60_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$388 U$$388/A1 U$$408/A2 U$$938/A1 U$$408/B2 VGND VGND VPWR VPWR U$$389/A sky130_fd_sc_hd__a22o_1
XU$$399 U$$399/A U$$411/A VGND VGND VPWR VPWR U$$399/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_24_clk _388_/CLK VGND VGND VPWR VPWR _382_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_79_5 dadda_fa_2_79_5/A dadda_fa_2_79_5/B dadda_fa_2_79_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_2/A dadda_fa_4_79_0/A sky130_fd_sc_hd__fa_2
XFILLER_113_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_2_30_4 U$$1663/X U$$1796/X VGND VGND VPWR VPWR dadda_fa_3_31_2/B dadda_fa_4_30_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_122_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_7_0_0 U$$7/X U$$9/B VGND VGND VPWR VPWR _297_/D _168_/D sky130_fd_sc_hd__ha_1
XFILLER_48_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1050 U$$1050/A U$$1094/B VGND VGND VPWR VPWR U$$1050/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_15_clk _370_/CLK VGND VGND VPWR VPWR _405_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1061 U$$924/A1 U$$1075/A2 U$$926/A1 U$$1075/B2 VGND VGND VPWR VPWR U$$1062/A sky130_fd_sc_hd__a22o_1
XU$$1072 U$$1072/A U$$962/A VGND VGND VPWR VPWR U$$1072/X sky130_fd_sc_hd__xor2_1
XU$$1083 U$$946/A1 U$$1093/A2 U$$948/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1084/A sky130_fd_sc_hd__a22o_1
XFILLER_149_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1094 U$$1094/A U$$1094/B VGND VGND VPWR VPWR U$$1094/X sky130_fd_sc_hd__xor2_1
XFILLER_164_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_82_7 U$$4028/X U$$4161/X VGND VGND VPWR VPWR dadda_fa_2_83_3/CIN dadda_fa_3_82_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_157_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_109_1 dadda_fa_5_109_1/A dadda_fa_5_109_1/B dadda_fa_5_109_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_110_0/B dadda_fa_7_109_0/A sky130_fd_sc_hd__fa_1
XFILLER_105_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_81_5 U$$3228/X U$$3361/X U$$3494/X VGND VGND VPWR VPWR dadda_fa_2_82_2/CIN
+ dadda_fa_2_81_5/B sky130_fd_sc_hd__fa_1
Xfanout602 U$$1785/X VGND VGND VPWR VPWR U$$1891/A2 sky130_fd_sc_hd__buf_6
XFILLER_132_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout613 U$$1593/A2 VGND VGND VPWR VPWR U$$1567/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout624 U$$141/X VGND VGND VPWR VPWR U$$259/A2 sky130_fd_sc_hd__buf_4
XFILLER_113_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout635 U$$1480/A2 VGND VGND VPWR VPWR U$$1502/A2 sky130_fd_sc_hd__buf_8
Xdadda_fa_1_74_4 U$$3347/X U$$3480/X U$$3613/X VGND VGND VPWR VPWR dadda_fa_2_75_1/CIN
+ dadda_fa_2_74_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_98_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout646 U$$1202/A2 VGND VGND VPWR VPWR U$$1194/A2 sky130_fd_sc_hd__buf_4
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout657 U$$1087/B2 VGND VGND VPWR VPWR U$$981/B2 sky130_fd_sc_hd__buf_6
Xfanout668 U$$807/B2 VGND VGND VPWR VPWR U$$763/B2 sky130_fd_sc_hd__buf_4
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_3 U$$3732/X U$$3865/X U$$3998/X VGND VGND VPWR VPWR dadda_fa_2_68_1/B
+ dadda_fa_2_67_4/B sky130_fd_sc_hd__fa_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout679 U$$553/X VGND VGND VPWR VPWR U$$676/B2 sky130_fd_sc_hd__buf_4
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_44_2 dadda_fa_4_44_2/A dadda_fa_4_44_2/B dadda_fa_4_44_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_45_0/CIN dadda_fa_5_44_1/CIN sky130_fd_sc_hd__fa_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_37_1 dadda_fa_4_37_1/A dadda_fa_4_37_1/B dadda_fa_4_37_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_38_0/B dadda_fa_5_37_1/B sky130_fd_sc_hd__fa_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_14_0 dadda_fa_7_14_0/A dadda_fa_7_14_0/B dadda_fa_7_14_0/CIN VGND VGND
+ VPWR VPWR _311_/D _182_/D sky130_fd_sc_hd__fa_1
XFILLER_27_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_270_ _408_/CLK _270_/D VGND VGND VPWR VPWR _270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_62_2 U$$929/X U$$1062/X U$$1195/X VGND VGND VPWR VPWR dadda_fa_1_63_6/A
+ dadda_fa_1_62_8/A sky130_fd_sc_hd__fa_1
XFILLER_49_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3903 U$$3903/A U$$3907/B VGND VGND VPWR VPWR U$$3903/X sky130_fd_sc_hd__xor2_1
XFILLER_76_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3914 U$$4462/A1 U$$3970/A2 U$$3916/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3915/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3925 U$$3925/A U$$3925/B VGND VGND VPWR VPWR U$$3925/X sky130_fd_sc_hd__xor2_1
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3936 U$$4484/A1 U$$3948/A2 U$$4484/B1 U$$3948/B2 VGND VGND VPWR VPWR U$$3937/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_32_0 U$$2269/B input182/X dadda_fa_3_32_0/CIN VGND VGND VPWR VPWR dadda_fa_4_33_0/B
+ dadda_fa_4_32_1/CIN sky130_fd_sc_hd__fa_1
XU$$3947 U$$3947/A U$$3949/B VGND VGND VPWR VPWR U$$3947/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$280 final_adder.U$$282/B final_adder.U$$280/B VGND VGND VPWR VPWR
+ final_adder.U$$406/B sky130_fd_sc_hd__and2_1
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3958 U$$4093/B1 U$$3960/A2 U$$3960/A1 U$$3960/B2 VGND VGND VPWR VPWR U$$3959/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$291 final_adder.U$$290/B final_adder.U$$165/X final_adder.U$$163/X
+ VGND VGND VPWR VPWR final_adder.U$$291/X sky130_fd_sc_hd__a21o_1
XU$$130 U$$539/B1 U$$98/A2 U$$406/A1 U$$98/B2 VGND VGND VPWR VPWR U$$131/A sky130_fd_sc_hd__a22o_1
XU$$3969 U$$3969/A U$$3972/A VGND VGND VPWR VPWR U$$3969/X sky130_fd_sc_hd__xor2_1
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$141 U$$139/Y U$$138/A U$$3/A U$$140/X U$$137/Y VGND VGND VPWR VPWR U$$141/X sky130_fd_sc_hd__a32o_4
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$152 U$$152/A U$$180/B VGND VGND VPWR VPWR U$$152/X sky130_fd_sc_hd__xor2_1
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$163 U$$26/A1 U$$213/A2 U$$28/A1 U$$213/B2 VGND VGND VPWR VPWR U$$164/A sky130_fd_sc_hd__a22o_1
XFILLER_73_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$174 U$$174/A U$$210/B VGND VGND VPWR VPWR U$$174/X sky130_fd_sc_hd__xor2_1
XFILLER_150_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$185 U$$868/B1 U$$219/A2 U$$735/A1 U$$219/B2 VGND VGND VPWR VPWR U$$186/A sky130_fd_sc_hd__a22o_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$196 U$$196/A U$$230/B VGND VGND VPWR VPWR U$$196/X sky130_fd_sc_hd__xor2_1
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_399_ _408_/CLK _399_/D VGND VGND VPWR VPWR _399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4395_1845 VGND VGND VPWR VPWR U$$4395_1845/HI U$$4395/B sky130_fd_sc_hd__conb_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_91_4 dadda_fa_2_91_4/A dadda_fa_2_91_4/B dadda_fa_2_91_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_92_1/CIN dadda_fa_3_91_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_84_3 dadda_fa_2_84_3/A dadda_fa_2_84_3/B dadda_fa_2_84_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_1/B dadda_fa_3_84_3/B sky130_fd_sc_hd__fa_1
Xdadda_fa_2_77_2 dadda_fa_2_77_2/A dadda_fa_2_77_2/B dadda_fa_2_77_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_1/A dadda_fa_3_77_3/A sky130_fd_sc_hd__fa_1
XFILLER_114_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_clk _201_/CLK VGND VGND VPWR VPWR _328_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_54_1 dadda_fa_5_54_1/A dadda_fa_5_54_1/B dadda_fa_5_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_55_0/B dadda_fa_7_54_0/A sky130_fd_sc_hd__fa_1
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_47_0 dadda_fa_5_47_0/A dadda_fa_5_47_0/B dadda_fa_5_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_48_0/A dadda_fa_6_47_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_100_1 U$$2867/X U$$3000/X U$$3133/X VGND VGND VPWR VPWR dadda_fa_3_101_1/CIN
+ dadda_fa_3_100_3/A sky130_fd_sc_hd__fa_1
XFILLER_24_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_121_0 U$$4372/X U$$4505/X input153/X VGND VGND VPWR VPWR dadda_fa_6_122_0/A
+ dadda_fa_6_121_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1408 U$$2739/A VGND VGND VPWR VPWR U$$2738/B sky130_fd_sc_hd__buf_6
Xfanout410 U$$676/A2 VGND VGND VPWR VPWR U$$674/A2 sky130_fd_sc_hd__buf_4
Xfanout1419 input31/X VGND VGND VPWR VPWR fanout1419/X sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_1_72_1 U$$2412/X U$$2545/X U$$2678/X VGND VGND VPWR VPWR dadda_fa_2_73_0/CIN
+ dadda_fa_2_72_3/CIN sky130_fd_sc_hd__fa_1
Xfanout421 U$$4369/A2 VGND VGND VPWR VPWR U$$4359/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout432 U$$415/X VGND VGND VPWR VPWR U$$545/A2 sky130_fd_sc_hd__buf_6
Xfanout443 U$$102/A2 VGND VGND VPWR VPWR U$$98/A2 sky130_fd_sc_hd__buf_4
XFILLER_24_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout454 U$$4057/A2 VGND VGND VPWR VPWR U$$4105/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_65_0 U$$2531/X U$$2664/X U$$2797/X VGND VGND VPWR VPWR dadda_fa_2_66_0/B
+ dadda_fa_2_65_3/B sky130_fd_sc_hd__fa_1
Xfanout465 U$$3966/A2 VGND VGND VPWR VPWR U$$3960/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout476 U$$3644/A2 VGND VGND VPWR VPWR U$$3604/A2 sky130_fd_sc_hd__buf_4
Xfanout487 U$$3429/X VGND VGND VPWR VPWR U$$3473/A2 sky130_fd_sc_hd__buf_4
XFILLER_86_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout498 U$$3422/A2 VGND VGND VPWR VPWR U$$3416/A2 sky130_fd_sc_hd__buf_4
XFILLER_171_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2509 U$$2509/A U$$2549/B VGND VGND VPWR VPWR U$$2509/X sky130_fd_sc_hd__xor2_1
XFILLER_73_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1808 U$$1808/A U$$1836/B VGND VGND VPWR VPWR U$$1808/X sky130_fd_sc_hd__xor2_1
XU$$1819 U$$997/A1 U$$1829/A2 U$$997/B1 U$$1829/B2 VGND VGND VPWR VPWR U$$1820/A sky130_fd_sc_hd__a22o_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_322_ _328_/CLK _322_/D VGND VGND VPWR VPWR _322_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_931 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_253_ _383_/CLK _253_/D VGND VGND VPWR VPWR _253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_184_ _321_/CLK _184_/D VGND VGND VPWR VPWR _184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_94_2 dadda_fa_3_94_2/A dadda_fa_3_94_2/B dadda_fa_3_94_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_1/A dadda_fa_4_94_2/B sky130_fd_sc_hd__fa_1
XFILLER_109_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_87_1 dadda_fa_3_87_1/A dadda_fa_3_87_1/B dadda_fa_3_87_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_0/CIN dadda_fa_4_87_2/A sky130_fd_sc_hd__fa_1
XFILLER_124_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_64_0 dadda_fa_6_64_0/A dadda_fa_6_64_0/B dadda_fa_6_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_65_0/B dadda_fa_7_64_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_9_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4401 U$$4401/A U$$4401/B VGND VGND VPWR VPWR U$$4401/X sky130_fd_sc_hd__xor2_1
XU$$4412 U$$4412/A1 U$$4388/X U$$4414/A1 U$$4458/B2 VGND VGND VPWR VPWR U$$4413/A
+ sky130_fd_sc_hd__a22o_1
XU$$4423 U$$4423/A U$$4423/B VGND VGND VPWR VPWR U$$4423/X sky130_fd_sc_hd__xor2_1
XU$$4434 U$$4434/A1 U$$4388/X U$$4436/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4435/A
+ sky130_fd_sc_hd__a22o_1
XU$$3700 input50/X VGND VGND VPWR VPWR U$$3702/B sky130_fd_sc_hd__inv_1
XFILLER_77_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4445 U$$4445/A U$$4445/B VGND VGND VPWR VPWR U$$4445/X sky130_fd_sc_hd__xor2_1
XFILLER_93_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3711 U$$3846/B1 U$$3791/A2 U$$3713/A1 U$$3791/B2 VGND VGND VPWR VPWR U$$3712/A
+ sky130_fd_sc_hd__a22o_1
XU$$4456 U$$4456/A1 U$$4388/X U$$4456/B1 U$$4389/X VGND VGND VPWR VPWR U$$4457/A sky130_fd_sc_hd__a22o_1
XU$$4467 U$$4467/A U$$4467/B VGND VGND VPWR VPWR U$$4467/X sky130_fd_sc_hd__xor2_1
XFILLER_37_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3722 U$$3722/A U$$3734/B VGND VGND VPWR VPWR U$$3722/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_116_1 U$$4229/X U$$4362/X U$$4495/X VGND VGND VPWR VPWR dadda_fa_5_117_0/B
+ dadda_fa_5_116_1/B sky130_fd_sc_hd__fa_1
XU$$3733 U$$3870/A1 U$$3757/A2 U$$3870/B1 U$$3757/B2 VGND VGND VPWR VPWR U$$3734/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4478 U$$4478/A1 U$$4388/X U$$4478/B1 U$$4488/B2 VGND VGND VPWR VPWR U$$4479/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_978 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3744 U$$3744/A U$$3790/B VGND VGND VPWR VPWR U$$3744/X sky130_fd_sc_hd__xor2_1
XFILLER_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4489 U$$4489/A U$$4489/B VGND VGND VPWR VPWR U$$4489/X sky130_fd_sc_hd__xor2_1
XU$$3755 U$$4027/B1 U$$3773/A2 U$$4440/B1 U$$3773/B2 VGND VGND VPWR VPWR U$$3756/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_109_0 dadda_fa_4_109_0/A dadda_fa_4_109_0/B dadda_fa_4_109_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_110_0/A dadda_fa_5_109_1/A sky130_fd_sc_hd__fa_1
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3766 U$$3766/A U$$3774/B VGND VGND VPWR VPWR U$$3766/X sky130_fd_sc_hd__xor2_1
XFILLER_33_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3777 U$$4462/A1 U$$3777/A2 U$$3916/A1 U$$3777/B2 VGND VGND VPWR VPWR U$$3778/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3788 U$$3788/A U$$3790/B VGND VGND VPWR VPWR U$$3788/X sky130_fd_sc_hd__xor2_1
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3799 U$$4482/B1 U$$3825/A2 U$$4349/A1 U$$3825/B2 VGND VGND VPWR VPWR U$$3800/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_82_0 U$$4294/X U$$4427/X input237/X VGND VGND VPWR VPWR dadda_fa_3_83_0/B
+ dadda_fa_3_82_2/B sky130_fd_sc_hd__fa_1
XFILLER_173_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_51_6 U$$2503/X U$$2636/X U$$2769/X VGND VGND VPWR VPWR dadda_fa_2_52_2/B
+ dadda_fa_2_51_5/B sky130_fd_sc_hd__fa_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_3_0 input190/X dadda_fa_7_3_0/B dadda_ha_6_3_0/SUM VGND VGND VPWR VPWR
+ _300_/D _171_/D sky130_fd_sc_hd__fa_1
XFILLER_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_81_0 dadda_fa_7_81_0/A dadda_fa_7_81_0/B dadda_fa_7_81_0/CIN VGND VGND
+ VPWR VPWR _378_/D _249_/D sky130_fd_sc_hd__fa_2
XFILLER_50_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_97_0 dadda_fa_4_97_0/A dadda_fa_4_97_0/B dadda_fa_4_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_98_0/A dadda_fa_5_97_1/A sky130_fd_sc_hd__fa_1
XFILLER_4_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1102_1782 VGND VGND VPWR VPWR U$$1102_1782/HI U$$1102/A1 sky130_fd_sc_hd__conb_1
XFILLER_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1205 input69/X VGND VGND VPWR VPWR U$$3870/A1 sky130_fd_sc_hd__buf_6
XFILLER_105_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1216 U$$4416/A1 VGND VGND VPWR VPWR U$$3181/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1227 U$$987/A1 VGND VGND VPWR VPWR U$$2631/A1 sky130_fd_sc_hd__buf_4
Xfanout1238 U$$8/A1 VGND VGND VPWR VPWR U$$965/B1 sky130_fd_sc_hd__buf_2
Xfanout1249 U$$651/B VGND VGND VPWR VPWR U$$639/B sky130_fd_sc_hd__buf_6
XFILLER_59_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3007 U$$3692/A1 U$$3011/A2 U$$3692/B1 U$$3011/B2 VGND VGND VPWR VPWR U$$3008/A
+ sky130_fd_sc_hd__a22o_1
XU$$3018 U$$3016/Y input39/X U$$3014/A U$$3017/X U$$3014/Y VGND VGND VPWR VPWR U$$3018/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3029 U$$3029/A U$$3061/B VGND VGND VPWR VPWR U$$3029/X sky130_fd_sc_hd__xor2_1
XFILLER_75_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2306 U$$2578/B1 U$$2310/A2 U$$2443/B1 U$$2310/B2 VGND VGND VPWR VPWR U$$2307/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2317 U$$2317/A U$$2328/A VGND VGND VPWR VPWR U$$2317/X sky130_fd_sc_hd__xor2_1
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2328 U$$2328/A VGND VGND VPWR VPWR U$$2328/Y sky130_fd_sc_hd__inv_1
XU$$2339 U$$3435/A1 U$$2413/A2 U$$971/A1 U$$2413/B2 VGND VGND VPWR VPWR U$$2340/A
+ sky130_fd_sc_hd__a22o_1
XU$$1605 U$$98/A1 U$$1641/A2 U$$98/B1 U$$1641/B2 VGND VGND VPWR VPWR U$$1606/A sky130_fd_sc_hd__a22o_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1616 U$$1616/A U$$1626/B VGND VGND VPWR VPWR U$$1616/X sky130_fd_sc_hd__xor2_1
XFILLER_43_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1627 U$$942/A1 U$$1635/A2 U$$2175/B1 U$$1635/B2 VGND VGND VPWR VPWR U$$1628/A
+ sky130_fd_sc_hd__a22o_1
XU$$1638 U$$1638/A U$$1644/A VGND VGND VPWR VPWR U$$1638/X sky130_fd_sc_hd__xor2_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1649 U$$1647/B U$$1630/B input17/X U$$1644/Y VGND VGND VPWR VPWR U$$1649/X sky130_fd_sc_hd__a22o_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_305_ _321_/CLK _305_/D VGND VGND VPWR VPWR _305_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_236_ _366_/CLK _236_/D VGND VGND VPWR VPWR _236_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_84_0_1925 VGND VGND VPWR VPWR dadda_fa_1_84_0/A dadda_fa_1_84_0_1925/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_971 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_61_5 dadda_fa_2_61_5/A dadda_fa_2_61_5/B dadda_fa_2_61_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_2/A dadda_fa_4_61_0/A sky130_fd_sc_hd__fa_2
XFILLER_66_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1750 U$$3382/B1 VGND VGND VPWR VPWR U$$4480/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_65_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_54_4 dadda_fa_2_54_4/A dadda_fa_2_54_4/B dadda_fa_2_54_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_1/CIN dadda_fa_3_54_3/CIN sky130_fd_sc_hd__fa_1
Xfanout1761 input102/X VGND VGND VPWR VPWR U$$914/B1 sky130_fd_sc_hd__buf_4
Xfanout1772 U$$3376/B1 VGND VGND VPWR VPWR U$$88/B1 sky130_fd_sc_hd__buf_4
XU$$4220 U$$4220/A1 U$$4236/A2 U$$4220/B1 U$$4236/B2 VGND VGND VPWR VPWR U$$4221/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4231 U$$4231/A U$$4231/B VGND VGND VPWR VPWR U$$4231/X sky130_fd_sc_hd__xor2_1
XU$$4242 U$$4377/B1 U$$4244/A2 U$$4244/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4243/A
+ sky130_fd_sc_hd__a22o_1
XU$$4253 U$$4253/A1 U$$4295/A2 U$$4392/A1 U$$4295/B2 VGND VGND VPWR VPWR U$$4254/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_47_3 dadda_fa_2_47_3/A dadda_fa_2_47_3/B dadda_fa_2_47_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_1/B dadda_fa_3_47_3/B sky130_fd_sc_hd__fa_1
XU$$4264 U$$4264/A U$$4292/B VGND VGND VPWR VPWR U$$4264/X sky130_fd_sc_hd__xor2_1
XU$$3530 U$$3530/A U$$3548/B VGND VGND VPWR VPWR U$$3530/X sky130_fd_sc_hd__xor2_1
XU$$4275 U$$4412/A1 U$$4325/A2 U$$4414/A1 U$$4325/B2 VGND VGND VPWR VPWR U$$4276/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4286 U$$4286/A U$$4383/A VGND VGND VPWR VPWR U$$4286/X sky130_fd_sc_hd__xor2_1
XU$$3541 U$$4226/A1 U$$3559/A2 U$$4226/B1 U$$3559/B2 VGND VGND VPWR VPWR U$$3542/A
+ sky130_fd_sc_hd__a22o_1
XU$$4297 U$$4434/A1 U$$4381/A2 U$$4436/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4298/A
+ sky130_fd_sc_hd__a22o_1
XU$$3552 U$$3552/A U$$3558/B VGND VGND VPWR VPWR U$$3552/X sky130_fd_sc_hd__xor2_1
XU$$3563 input48/X VGND VGND VPWR VPWR U$$3565/B sky130_fd_sc_hd__inv_1
XFILLER_80_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3574 U$$3846/B1 U$$3658/A2 U$$3713/A1 U$$3658/B2 VGND VGND VPWR VPWR U$$3575/A
+ sky130_fd_sc_hd__a22o_1
XU$$1641_1791 VGND VGND VPWR VPWR U$$1641_1791/HI U$$1641/B1 sky130_fd_sc_hd__conb_1
XU$$2840 U$$2840/A1 U$$2840/A2 U$$2840/B1 U$$2840/B2 VGND VGND VPWR VPWR U$$2841/A
+ sky130_fd_sc_hd__a22o_1
XU$$3585 U$$3585/A U$$3601/B VGND VGND VPWR VPWR U$$3585/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_17_1 dadda_fa_5_17_1/A dadda_fa_5_17_1/B dadda_fa_5_17_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_18_0/B dadda_fa_7_17_0/A sky130_fd_sc_hd__fa_1
XU$$3596 U$$3870/A1 U$$3604/A2 U$$3870/B1 U$$3604/B2 VGND VGND VPWR VPWR U$$3597/A
+ sky130_fd_sc_hd__a22o_1
XU$$2851 U$$2851/A U$$2876/A VGND VGND VPWR VPWR U$$2851/X sky130_fd_sc_hd__xor2_1
XU$$2862 U$$3684/A1 U$$2872/A2 U$$2862/B1 U$$2872/B2 VGND VGND VPWR VPWR U$$2863/A
+ sky130_fd_sc_hd__a22o_1
XU$$2873 U$$2873/A U$$2873/B VGND VGND VPWR VPWR U$$2873/X sky130_fd_sc_hd__xor2_1
XU$$2884 U$$2884/A U$$2926/B VGND VGND VPWR VPWR U$$2884/X sky130_fd_sc_hd__xor2_1
XU$$2895 U$$3030/B1 U$$2929/A2 U$$2897/A1 U$$2929/B2 VGND VGND VPWR VPWR U$$2896/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_4_120_1 U$$4237/X U$$4370/X VGND VGND VPWR VPWR dadda_fa_5_121_1/B dadda_ha_4_120_1/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_103_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_43_4 U$$1689/X U$$1822/X VGND VGND VPWR VPWR dadda_fa_2_44_4/A dadda_fa_3_43_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_88_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$813 final_adder.U$$780/A final_adder.U$$733/X final_adder.U$$701/X
+ VGND VGND VPWR VPWR final_adder.U$$813/X sky130_fd_sc_hd__a21o_1
XFILLER_21_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_4_13_2 U$$831/X input161/X VGND VGND VPWR VPWR dadda_fa_5_14_0/CIN dadda_ha_4_13_2/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_56_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$857 final_adder.U$$760/X final_adder.U$$825/X final_adder.U$$761/X
+ VGND VGND VPWR VPWR final_adder.U$$857/X sky130_fd_sc_hd__a21o_1
XFILLER_57_978 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$707 U$$707/A1 U$$771/A2 U$$709/A1 U$$771/B2 VGND VGND VPWR VPWR U$$708/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$879 final_adder.U$$782/X final_adder.U$$735/X final_adder.U$$783/X
+ VGND VGND VPWR VPWR final_adder.U$$879/X sky130_fd_sc_hd__a21o_1
XU$$718 U$$718/A U$$764/B VGND VGND VPWR VPWR U$$718/X sky130_fd_sc_hd__xor2_1
XU$$729 U$$864/B1 U$$763/A2 U$$729/B1 U$$763/B2 VGND VGND VPWR VPWR U$$730/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_42_2 U$$889/X U$$1022/X U$$1155/X VGND VGND VPWR VPWR dadda_fa_2_43_3/CIN
+ dadda_fa_2_42_5/B sky130_fd_sc_hd__fa_1
XFILLER_83_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_12_0 U$$31/X U$$164/X U$$297/X VGND VGND VPWR VPWR dadda_fa_5_13_0/A dadda_fa_5_12_1/A
+ sky130_fd_sc_hd__fa_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_72_0_1920 VGND VGND VPWR VPWR dadda_fa_0_72_0/A dadda_fa_0_72_0_1920/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1002 input92/X VGND VGND VPWR VPWR fanout999/A sky130_fd_sc_hd__buf_8
Xdadda_fa_3_64_3 dadda_fa_3_64_3/A dadda_fa_3_64_3/B dadda_fa_3_64_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_1/B dadda_fa_4_64_2/CIN sky130_fd_sc_hd__fa_1
Xfanout1013 U$$4182/A1 VGND VGND VPWR VPWR U$$70/B1 sky130_fd_sc_hd__buf_6
XFILLER_79_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1024 input9/X VGND VGND VPWR VPWR U$$1189/B sky130_fd_sc_hd__buf_4
XFILLER_120_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1035 U$$4315/B1 VGND VGND VPWR VPWR U$$4454/A1 sky130_fd_sc_hd__buf_4
Xfanout1046 U$$4257/B1 VGND VGND VPWR VPWR U$$3163/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1057 U$$3080/A1 VGND VGND VPWR VPWR U$$612/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_57_2 dadda_fa_3_57_2/A dadda_fa_3_57_2/B dadda_fa_3_57_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_1/A dadda_fa_4_57_2/B sky130_fd_sc_hd__fa_1
XFILLER_0_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1068 U$$4446/B1 VGND VGND VPWR VPWR U$$4174/A1 sky130_fd_sc_hd__buf_2
XFILLER_86_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1079 U$$3072/B1 VGND VGND VPWR VPWR U$$469/B1 sky130_fd_sc_hd__buf_4
XFILLER_75_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_27_0 dadda_fa_6_27_0/A dadda_fa_6_27_0/B dadda_fa_6_27_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_28_0/B dadda_fa_7_27_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2103 U$$870/A1 U$$2107/A2 U$$872/A1 U$$2107/B2 VGND VGND VPWR VPWR U$$2104/A sky130_fd_sc_hd__a22o_1
XFILLER_63_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2114 U$$2114/A U$$2148/B VGND VGND VPWR VPWR U$$2114/X sky130_fd_sc_hd__xor2_1
XFILLER_34_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2125 U$$70/A1 U$$2139/A2 U$$70/B1 U$$2139/B2 VGND VGND VPWR VPWR U$$2126/A sky130_fd_sc_hd__a22o_1
XU$$2136 U$$2136/A U$$2140/B VGND VGND VPWR VPWR U$$2136/X sky130_fd_sc_hd__xor2_1
XU$$1402 U$$443/A1 U$$1414/A2 U$$34/A1 U$$1414/B2 VGND VGND VPWR VPWR U$$1403/A sky130_fd_sc_hd__a22o_1
XU$$2147 U$$640/A1 U$$2147/A2 U$$916/A1 U$$2147/B2 VGND VGND VPWR VPWR U$$2148/A sky130_fd_sc_hd__a22o_1
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2158 U$$2158/A U$$2191/A VGND VGND VPWR VPWR U$$2158/X sky130_fd_sc_hd__xor2_1
XU$$1413 U$$1413/A U$$1415/B VGND VGND VPWR VPWR U$$1413/X sky130_fd_sc_hd__xor2_1
XU$$1424 U$$465/A1 U$$1426/A2 U$$465/B1 U$$1426/B2 VGND VGND VPWR VPWR U$$1425/A sky130_fd_sc_hd__a22o_1
XFILLER_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2169 U$$388/A1 U$$2177/A2 U$$2443/B1 U$$2177/B2 VGND VGND VPWR VPWR U$$2170/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1435 U$$1435/A U$$1461/B VGND VGND VPWR VPWR U$$1435/X sky130_fd_sc_hd__xor2_1
XU$$1446 U$$76/A1 U$$1480/A2 U$$78/A1 U$$1480/B2 VGND VGND VPWR VPWR U$$1447/A sky130_fd_sc_hd__a22o_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1457 U$$1457/A U$$1461/B VGND VGND VPWR VPWR U$$1457/X sky130_fd_sc_hd__xor2_1
XU$$1468 U$$98/A1 U$$1504/A2 U$$98/B1 U$$1504/B2 VGND VGND VPWR VPWR U$$1469/A sky130_fd_sc_hd__a22o_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1479 U$$1479/A U$$1491/B VGND VGND VPWR VPWR U$$1479/X sky130_fd_sc_hd__xor2_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_219_ _348_/CLK _219_/D VGND VGND VPWR VPWR _219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$109 _405_/Q _277_/Q VGND VGND VPWR VPWR final_adder.U$$147/B1 final_adder.U$$146/B
+ sky130_fd_sc_hd__ha_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_52_1 dadda_fa_2_52_1/A dadda_fa_2_52_1/B dadda_fa_2_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_0/CIN dadda_fa_3_52_2/CIN sky130_fd_sc_hd__fa_1
Xfanout1580 U$$3580/A1 VGND VGND VPWR VPWR U$$840/A1 sky130_fd_sc_hd__buf_4
Xfanout1591 input12/X VGND VGND VPWR VPWR U$$121/B sky130_fd_sc_hd__buf_8
XU$$4050 U$$4050/A U$$4098/B VGND VGND VPWR VPWR U$$4050/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_45_0 U$$2358/X U$$2491/X U$$2624/X VGND VGND VPWR VPWR dadda_fa_3_46_0/B
+ dadda_fa_3_45_2/B sky130_fd_sc_hd__fa_1
XFILLER_39_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4061 U$$4196/B1 U$$4081/A2 U$$4198/B1 U$$4081/B2 VGND VGND VPWR VPWR U$$4062/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4072 U$$4072/A U$$4094/B VGND VGND VPWR VPWR U$$4072/X sky130_fd_sc_hd__xor2_1
XU$$4083 U$$4220/A1 U$$4105/A2 U$$4220/B1 U$$4105/B2 VGND VGND VPWR VPWR U$$4084/A
+ sky130_fd_sc_hd__a22o_1
XU$$4094 U$$4094/A U$$4094/B VGND VGND VPWR VPWR U$$4094/X sky130_fd_sc_hd__xor2_1
XU$$3360 U$$3495/B1 U$$3372/A2 U$$3499/A1 U$$3372/B2 VGND VGND VPWR VPWR U$$3361/A
+ sky130_fd_sc_hd__a22o_1
XU$$3371 U$$3371/A U$$3373/B VGND VGND VPWR VPWR U$$3371/X sky130_fd_sc_hd__xor2_1
XU$$3382 U$$3382/A1 U$$3422/A2 U$$3382/B1 U$$3422/B2 VGND VGND VPWR VPWR U$$3383/A
+ sky130_fd_sc_hd__a22o_1
XU$$3393 U$$3393/A U$$3417/B VGND VGND VPWR VPWR U$$3393/X sky130_fd_sc_hd__xor2_1
XFILLER_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2670 U$$2670/A U$$2740/A VGND VGND VPWR VPWR U$$2670/X sky130_fd_sc_hd__xor2_1
XFILLER_62_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2681 U$$215/A1 U$$2681/A2 U$$80/A1 U$$2681/B2 VGND VGND VPWR VPWR U$$2682/A sky130_fd_sc_hd__a22o_1
XU$$2692 U$$2692/A U$$2740/A VGND VGND VPWR VPWR U$$2692/X sky130_fd_sc_hd__xor2_1
XU$$1980 U$$882/B1 U$$1980/A2 U$$747/B1 U$$1980/B2 VGND VGND VPWR VPWR U$$1981/A sky130_fd_sc_hd__a22o_1
XFILLER_21_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1991 U$$1991/A U$$2007/B VGND VGND VPWR VPWR U$$1991/X sky130_fd_sc_hd__xor2_1
XFILLER_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2737_1808 VGND VGND VPWR VPWR U$$2737_1808/HI U$$2737/B1 sky130_fd_sc_hd__conb_1
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_74_2 dadda_fa_4_74_2/A dadda_fa_4_74_2/B dadda_fa_4_74_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_75_0/CIN dadda_fa_5_74_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_67_1 dadda_fa_4_67_1/A dadda_fa_4_67_1/B dadda_fa_4_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_68_0/B dadda_fa_5_67_1/B sky130_fd_sc_hd__fa_1
XFILLER_131_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput105 b[46] VGND VGND VPWR VPWR input105/X sky130_fd_sc_hd__buf_6
Xinput116 b[56] VGND VGND VPWR VPWR input116/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_7_44_0 dadda_fa_7_44_0/A dadda_fa_7_44_0/B dadda_fa_7_44_0/CIN VGND VGND
+ VPWR VPWR _341_/D _212_/D sky130_fd_sc_hd__fa_1
XFILLER_89_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput127 b[8] VGND VGND VPWR VPWR input127/X sky130_fd_sc_hd__buf_2
Xinput138 c[108] VGND VGND VPWR VPWR input138/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_34_0 U$$75/X U$$208/X VGND VGND VPWR VPWR dadda_fa_2_35_5/CIN dadda_fa_3_34_0/A
+ sky130_fd_sc_hd__ha_1
Xinput149 c[118] VGND VGND VPWR VPWR input149/X sky130_fd_sc_hd__buf_2
XFILLER_102_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$610 final_adder.U$$610/A final_adder.U$$610/B VGND VGND VPWR VPWR
+ final_adder.U$$714/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$621 final_adder.U$$612/A final_adder.U$$505/X final_adder.U$$497/X
+ VGND VGND VPWR VPWR final_adder.U$$621/X sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$632 final_adder.U$$648/B final_adder.U$$632/B VGND VGND VPWR VPWR
+ final_adder.U$$744/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$643 final_adder.U$$642/B final_adder.U$$539/X final_adder.U$$523/X
+ VGND VGND VPWR VPWR final_adder.U$$643/X sky130_fd_sc_hd__a21o_1
XFILLER_56_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$654 final_adder.U$$670/B final_adder.U$$654/B VGND VGND VPWR VPWR
+ final_adder.U$$766/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$665 final_adder.U$$664/B final_adder.U$$561/X final_adder.U$$545/X
+ VGND VGND VPWR VPWR final_adder.U$$665/X sky130_fd_sc_hd__a21o_1
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$504 U$$504/A U$$504/B VGND VGND VPWR VPWR U$$504/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$676 final_adder.U$$692/B final_adder.U$$676/B VGND VGND VPWR VPWR
+ final_adder.U$$788/B sky130_fd_sc_hd__and2_1
XU$$515 U$$650/B1 U$$545/A2 U$$517/A1 U$$545/B2 VGND VGND VPWR VPWR U$$516/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$687 final_adder.U$$686/B final_adder.U$$583/X final_adder.U$$567/X
+ VGND VGND VPWR VPWR final_adder.U$$687/X sky130_fd_sc_hd__a21o_1
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$526 U$$526/A U$$536/B VGND VGND VPWR VPWR U$$526/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$698 final_adder.U$$714/B final_adder.U$$698/B VGND VGND VPWR VPWR
+ final_adder.U$$778/A sky130_fd_sc_hd__and2_1
XU$$537 U$$672/B1 U$$539/A2 U$$539/A1 U$$539/B2 VGND VGND VPWR VPWR U$$538/A sky130_fd_sc_hd__a22o_1
XFILLER_72_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$548 U$$548/A VGND VGND VPWR VPWR U$$548/Y sky130_fd_sc_hd__inv_1
XU$$559 U$$559/A U$$607/B VGND VGND VPWR VPWR U$$559/X sky130_fd_sc_hd__xor2_1
XFILLER_13_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_62_0 dadda_fa_3_62_0/A dadda_fa_3_62_0/B dadda_fa_3_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_0/B dadda_fa_4_62_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_859 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_4_9_0 U$$25/X U$$158/X VGND VGND VPWR VPWR dadda_fa_5_10_1/A dadda_ha_4_9_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$1210 U$$386/B1 U$$1226/A2 U$$253/A1 U$$1226/B2 VGND VGND VPWR VPWR U$$1211/A sky130_fd_sc_hd__a22o_1
XFILLER_90_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1221 U$$1221/A U$$1221/B VGND VGND VPWR VPWR U$$1221/X sky130_fd_sc_hd__xor2_1
XU$$1232 U$$1233/A VGND VGND VPWR VPWR U$$1232/Y sky130_fd_sc_hd__inv_1
XU$$1243 U$$3435/A1 U$$1309/A2 U$$697/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1244/A
+ sky130_fd_sc_hd__a22o_1
XU$$1254 U$$1254/A U$$1300/B VGND VGND VPWR VPWR U$$1254/X sky130_fd_sc_hd__xor2_1
XU$$1265 U$$991/A1 U$$1295/A2 U$$993/A1 U$$1295/B2 VGND VGND VPWR VPWR U$$1266/A sky130_fd_sc_hd__a22o_1
XU$$1276 U$$1276/A U$$1278/B VGND VGND VPWR VPWR U$$1276/X sky130_fd_sc_hd__xor2_1
XU$$1287 U$$465/A1 U$$1295/A2 U$$465/B1 U$$1295/B2 VGND VGND VPWR VPWR U$$1288/A sky130_fd_sc_hd__a22o_1
XU$$1298 U$$1298/A U$$1328/B VGND VGND VPWR VPWR U$$1298/X sky130_fd_sc_hd__xor2_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1376_1787 VGND VGND VPWR VPWR U$$1376_1787/HI U$$1376/A1 sky130_fd_sc_hd__conb_1
Xdadda_fa_5_84_1 dadda_fa_5_84_1/A dadda_fa_5_84_1/B dadda_fa_5_84_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_85_0/B dadda_fa_7_84_0/A sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$1070 final_adder.U$$208/A final_adder.U$$821/X VGND VGND VPWR VPWR
+ output325/A sky130_fd_sc_hd__xor2_1
XFILLER_116_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1081 final_adder.U$$198/B final_adder.U$$969/X VGND VGND VPWR VPWR
+ output337/A sky130_fd_sc_hd__xor2_1
XFILLER_117_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1092 final_adder.U$$186/A final_adder.U$$895/X VGND VGND VPWR VPWR
+ output349/A sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_77_0 dadda_fa_5_77_0/A dadda_fa_5_77_0/B dadda_fa_5_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_78_0/A dadda_fa_6_77_0/CIN sky130_fd_sc_hd__fa_1
Xfanout806 U$$2608/X VGND VGND VPWR VPWR U$$2707/B2 sky130_fd_sc_hd__buf_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout817 fanout820/X VGND VGND VPWR VPWR U$$2548/B2 sky130_fd_sc_hd__clkbuf_4
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout828 U$$2334/X VGND VGND VPWR VPWR U$$2463/B2 sky130_fd_sc_hd__buf_6
XFILLER_97_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_76_8 dadda_fa_1_76_8/A dadda_fa_1_76_8/B dadda_fa_1_76_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_77_3/A dadda_fa_3_76_0/A sky130_fd_sc_hd__fa_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout839 U$$2147/B2 VGND VGND VPWR VPWR U$$2107/B2 sky130_fd_sc_hd__buf_6
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_7 dadda_fa_1_69_7/A dadda_fa_1_69_7/B dadda_fa_1_69_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_70_2/CIN dadda_fa_2_69_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3190 U$$3190/A U$$3196/B VGND VGND VPWR VPWR U$$3190/X sky130_fd_sc_hd__xor2_1
XFILLER_41_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2600_1805 VGND VGND VPWR VPWR U$$2600_1805/HI U$$2600/B1 sky130_fd_sc_hd__conb_1
XFILLER_148_894 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_100_3 dadda_fa_3_100_3/A dadda_fa_3_100_3/B dadda_fa_3_100_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_101_1/B dadda_fa_4_100_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_95_0 U$$2191/Y U$$2325/X U$$2458/X VGND VGND VPWR VPWR dadda_fa_2_96_5/CIN
+ dadda_fa_3_95_0/A sky130_fd_sc_hd__fa_1
XFILLER_174_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_2_108_0 dadda_ha_2_108_0/A U$$3149/X VGND VGND VPWR VPWR dadda_fa_4_109_0/A
+ dadda_fa_4_108_0/A sky130_fd_sc_hd__ha_1
XFILLER_76_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$440 final_adder.U$$444/B final_adder.U$$440/B VGND VGND VPWR VPWR
+ final_adder.U$$564/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$451 final_adder.U$$450/B final_adder.U$$329/X final_adder.U$$325/X
+ VGND VGND VPWR VPWR final_adder.U$$451/X sky130_fd_sc_hd__a21o_1
XFILLER_29_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$462 final_adder.U$$466/B final_adder.U$$462/B VGND VGND VPWR VPWR
+ final_adder.U$$586/B sky130_fd_sc_hd__and2_1
XFILLER_18_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$301 U$$301/A U$$341/B VGND VGND VPWR VPWR U$$301/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_107_0 dadda_fa_6_107_0/A dadda_fa_6_107_0/B dadda_fa_6_107_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_108_0/B dadda_fa_7_107_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$473 final_adder.U$$472/B final_adder.U$$351/X final_adder.U$$347/X
+ VGND VGND VPWR VPWR final_adder.U$$473/X sky130_fd_sc_hd__a21o_1
XFILLER_45_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$312 U$$447/B1 U$$312/A2 U$$314/A1 U$$312/B2 VGND VGND VPWR VPWR U$$313/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$484 final_adder.U$$488/B final_adder.U$$484/B VGND VGND VPWR VPWR
+ final_adder.U$$608/B sky130_fd_sc_hd__and2_1
XFILLER_17_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$323 U$$323/A U$$353/B VGND VGND VPWR VPWR U$$323/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$495 final_adder.U$$494/B final_adder.U$$373/X final_adder.U$$369/X
+ VGND VGND VPWR VPWR final_adder.U$$495/X sky130_fd_sc_hd__a21o_1
XU$$334 U$$469/B1 U$$352/A2 U$$884/A1 U$$352/B2 VGND VGND VPWR VPWR U$$335/A sky130_fd_sc_hd__a22o_1
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$345 U$$345/A U$$347/B VGND VGND VPWR VPWR U$$345/X sky130_fd_sc_hd__xor2_1
XU$$356 U$$765/B1 U$$362/A2 U$$632/A1 U$$362/B2 VGND VGND VPWR VPWR U$$357/A sky130_fd_sc_hd__a22o_1
XFILLER_33_918 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_27_3 dadda_fa_3_27_3/A dadda_fa_3_27_3/B dadda_fa_3_27_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_28_1/B dadda_fa_4_27_2/CIN sky130_fd_sc_hd__fa_1
XU$$367 U$$367/A U$$407/B VGND VGND VPWR VPWR U$$367/X sky130_fd_sc_hd__xor2_1
XU$$378 U$$650/B1 U$$386/A2 U$$517/A1 U$$386/B2 VGND VGND VPWR VPWR U$$379/A sky130_fd_sc_hd__a22o_1
XFILLER_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$389 U$$389/A U$$410/A VGND VGND VPWR VPWR U$$389/X sky130_fd_sc_hd__xor2_1
XFILLER_60_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_94_0 dadda_fa_6_94_0/A dadda_fa_6_94_0/B dadda_fa_6_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_95_0/B dadda_fa_7_94_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_145_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$890 U$$66/B1 U$$898/A2 U$$892/A1 U$$898/B2 VGND VGND VPWR VPWR U$$891/A sky130_fd_sc_hd__a22o_1
XU$$1040 U$$1040/A U$$1046/B VGND VGND VPWR VPWR U$$1040/X sky130_fd_sc_hd__xor2_1
XU$$1051 U$$640/A1 U$$1093/A2 U$$916/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1052/A sky130_fd_sc_hd__a22o_1
XU$$1062 U$$1062/A U$$1062/B VGND VGND VPWR VPWR U$$1062/X sky130_fd_sc_hd__xor2_1
XU$$1073 U$$388/A1 U$$1075/A2 U$$936/B1 U$$1075/B2 VGND VGND VPWR VPWR U$$1074/A sky130_fd_sc_hd__a22o_1
XU$$1084 U$$1084/A U$$1094/B VGND VGND VPWR VPWR U$$1084/X sky130_fd_sc_hd__xor2_1
XU$$1095 U$$990/B VGND VGND VPWR VPWR U$$1095/Y sky130_fd_sc_hd__inv_1
XFILLER_149_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_81_6 U$$3627/X U$$3760/X U$$3893/X VGND VGND VPWR VPWR dadda_fa_2_82_3/A
+ dadda_fa_2_81_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout603 U$$1726/A2 VGND VGND VPWR VPWR U$$1696/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout614 U$$1621/A2 VGND VGND VPWR VPWR U$$1593/A2 sky130_fd_sc_hd__buf_2
XFILLER_99_973 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_74_5 U$$3746/X U$$3879/X U$$4012/X VGND VGND VPWR VPWR dadda_fa_2_75_2/A
+ dadda_fa_2_74_5/A sky130_fd_sc_hd__fa_1
Xfanout625 U$$213/A2 VGND VGND VPWR VPWR U$$179/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout636 U$$1374/X VGND VGND VPWR VPWR U$$1480/A2 sky130_fd_sc_hd__buf_8
XFILLER_113_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout647 U$$1202/A2 VGND VGND VPWR VPWR U$$1230/A2 sky130_fd_sc_hd__buf_6
Xfanout658 U$$1087/B2 VGND VGND VPWR VPWR U$$1093/B2 sky130_fd_sc_hd__buf_6
XU$$4413_1854 VGND VGND VPWR VPWR U$$4413_1854/HI U$$4413/B sky130_fd_sc_hd__conb_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_4 U$$4131/X U$$4264/X U$$4397/X VGND VGND VPWR VPWR dadda_fa_2_68_1/CIN
+ dadda_fa_2_67_4/CIN sky130_fd_sc_hd__fa_1
Xfanout669 U$$807/B2 VGND VGND VPWR VPWR U$$769/B2 sky130_fd_sc_hd__buf_4
XFILLER_86_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_37_2 dadda_fa_4_37_2/A dadda_fa_4_37_2/B dadda_fa_4_37_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_38_0/CIN dadda_fa_5_37_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_0_63_5 U$$2128/X U$$2261/X VGND VGND VPWR VPWR dadda_fa_1_64_7/A dadda_fa_2_63_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_150_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_62_3 U$$1328/X U$$1461/X U$$1594/X VGND VGND VPWR VPWR dadda_fa_1_63_6/B
+ dadda_fa_1_62_8/B sky130_fd_sc_hd__fa_1
XFILLER_37_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3904 U$$4176/B1 U$$3906/A2 U$$4043/A1 U$$3906/B2 VGND VGND VPWR VPWR U$$3905/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3915 U$$3915/A U$$3965/B VGND VGND VPWR VPWR U$$3915/X sky130_fd_sc_hd__xor2_1
XU$$3926 U$$4198/B1 U$$3948/A2 U$$4476/A1 U$$3948/B2 VGND VGND VPWR VPWR U$$3927/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3937 U$$3937/A U$$3949/B VGND VGND VPWR VPWR U$$3937/X sky130_fd_sc_hd__xor2_1
XFILLER_18_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$270 final_adder.U$$272/B final_adder.U$$270/B VGND VGND VPWR VPWR
+ final_adder.U$$396/B sky130_fd_sc_hd__and2_1
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3948 U$$3948/A1 U$$3948/A2 U$$3948/B1 U$$3948/B2 VGND VGND VPWR VPWR U$$3949/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$281 final_adder.U$$280/B final_adder.U$$155/X final_adder.U$$153/X
+ VGND VGND VPWR VPWR final_adder.U$$281/X sky130_fd_sc_hd__a21o_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_32_1 dadda_fa_3_32_1/A dadda_fa_3_32_1/B dadda_fa_3_32_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_33_0/CIN dadda_fa_4_32_2/A sky130_fd_sc_hd__fa_2
XU$$120 U$$120/A1 U$$120/A2 U$$120/B1 U$$120/B2 VGND VGND VPWR VPWR U$$121/A sky130_fd_sc_hd__a22o_1
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$292 final_adder.U$$294/B final_adder.U$$292/B VGND VGND VPWR VPWR
+ final_adder.U$$418/B sky130_fd_sc_hd__and2_1
XU$$131 U$$131/A U$$3/A VGND VGND VPWR VPWR U$$131/X sky130_fd_sc_hd__xor2_1
XU$$3959 U$$3959/A U$$3961/B VGND VGND VPWR VPWR U$$3959/X sky130_fd_sc_hd__xor2_1
XU$$142 U$$140/B U$$3/A U$$138/A U$$137/Y VGND VGND VPWR VPWR U$$142/X sky130_fd_sc_hd__a22o_2
XFILLER_73_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$153 U$$16/A1 U$$179/A2 U$$18/A1 U$$179/B2 VGND VGND VPWR VPWR U$$154/A sky130_fd_sc_hd__a22o_1
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_25_0 U$$722/X U$$855/X U$$988/X VGND VGND VPWR VPWR dadda_fa_4_26_0/B
+ dadda_fa_4_25_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$164 U$$164/A U$$214/B VGND VGND VPWR VPWR U$$164/X sky130_fd_sc_hd__xor2_1
XFILLER_72_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$175 U$$447/B1 U$$207/A2 U$$314/A1 U$$207/B2 VGND VGND VPWR VPWR U$$176/A sky130_fd_sc_hd__a22o_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$186 U$$186/A U$$220/B VGND VGND VPWR VPWR U$$186/X sky130_fd_sc_hd__xor2_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$197 U$$60/A1 U$$229/A2 U$$62/A1 U$$229/B2 VGND VGND VPWR VPWR U$$198/A sky130_fd_sc_hd__a22o_1
XFILLER_72_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_398_ _408_/CLK _398_/D VGND VGND VPWR VPWR _398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_120_0_1940 VGND VGND VPWR VPWR dadda_fa_4_120_0/A dadda_fa_4_120_0_1940/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_126_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_91_5 dadda_fa_2_91_5/A dadda_fa_2_91_5/B dadda_fa_2_91_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_92_2/A dadda_fa_4_91_0/A sky130_fd_sc_hd__fa_1
XFILLER_5_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_84_4 dadda_fa_2_84_4/A dadda_fa_2_84_4/B dadda_fa_2_84_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_1/CIN dadda_fa_3_84_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_126_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_77_3 dadda_fa_2_77_3/A dadda_fa_2_77_3/B dadda_fa_2_77_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_1/B dadda_fa_3_77_3/B sky130_fd_sc_hd__fa_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_47_1 dadda_fa_5_47_1/A dadda_fa_5_47_1/B dadda_fa_5_47_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_48_0/B dadda_fa_7_47_0/A sky130_fd_sc_hd__fa_1
XFILLER_110_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_100_2 U$$3266/X U$$3399/X U$$3532/X VGND VGND VPWR VPWR dadda_fa_3_101_2/A
+ dadda_fa_3_100_3/B sky130_fd_sc_hd__fa_1
XFILLER_51_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4443_1869 VGND VGND VPWR VPWR U$$4443_1869/HI U$$4443/B sky130_fd_sc_hd__conb_1
XFILLER_32_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_121_1 dadda_fa_5_121_1/A dadda_fa_5_121_1/B dadda_fa_5_121_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_122_0/B dadda_fa_7_121_0/A sky130_fd_sc_hd__fa_1
XFILLER_139_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_114_0 dadda_fa_5_114_0/A dadda_fa_5_114_0/B dadda_fa_5_114_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_115_0/A dadda_fa_6_114_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_164_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout400 U$$807/A2 VGND VGND VPWR VPWR U$$763/A2 sky130_fd_sc_hd__buf_4
Xfanout411 U$$552/X VGND VGND VPWR VPWR U$$676/A2 sky130_fd_sc_hd__buf_4
Xfanout1409 U$$2745/A2 VGND VGND VPWR VPWR U$$2739/A sky130_fd_sc_hd__buf_6
Xfanout422 U$$4325/A2 VGND VGND VPWR VPWR U$$4369/A2 sky130_fd_sc_hd__buf_2
XFILLER_132_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_72_2 U$$2811/X U$$2944/X U$$3077/X VGND VGND VPWR VPWR dadda_fa_2_73_1/A
+ dadda_fa_2_72_4/A sky130_fd_sc_hd__fa_1
Xfanout433 U$$4244/A2 VGND VGND VPWR VPWR U$$4158/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_132_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout444 U$$48/A2 VGND VGND VPWR VPWR U$$8/A2 sky130_fd_sc_hd__buf_2
Xfanout455 U$$3977/X VGND VGND VPWR VPWR U$$4107/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_65_1 U$$2930/X U$$3063/X U$$3196/X VGND VGND VPWR VPWR dadda_fa_2_66_0/CIN
+ dadda_fa_2_65_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout466 U$$3924/A2 VGND VGND VPWR VPWR U$$3966/A2 sky130_fd_sc_hd__buf_2
Xfanout477 U$$3644/A2 VGND VGND VPWR VPWR U$$3640/A2 sky130_fd_sc_hd__buf_4
XFILLER_101_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout488 U$$3439/A2 VGND VGND VPWR VPWR U$$3523/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_4_42_0 dadda_fa_4_42_0/A dadda_fa_4_42_0/B dadda_fa_4_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_43_0/A dadda_fa_5_42_1/A sky130_fd_sc_hd__fa_1
Xfanout499 U$$3422/A2 VGND VGND VPWR VPWR U$$3418/A2 sky130_fd_sc_hd__buf_2
Xdadda_fa_1_58_0 U$$1586/X U$$1719/X U$$1852/X VGND VGND VPWR VPWR dadda_fa_2_59_0/B
+ dadda_fa_2_58_3/B sky130_fd_sc_hd__fa_1
XFILLER_58_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1809 U$$576/A1 U$$1881/A2 U$$576/B1 U$$1881/B2 VGND VGND VPWR VPWR U$$1810/A sky130_fd_sc_hd__a22o_1
XFILLER_54_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_321_ _321_/CLK _321_/D VGND VGND VPWR VPWR _321_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_252_ _380_/CLK _252_/D VGND VGND VPWR VPWR _252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_183_ _328_/CLK _183_/D VGND VGND VPWR VPWR _183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_94_3 dadda_fa_3_94_3/A dadda_fa_3_94_3/B dadda_fa_3_94_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_1/B dadda_fa_4_94_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_109_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_87_2 dadda_fa_3_87_2/A dadda_fa_3_87_2/B dadda_fa_3_87_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_1/A dadda_fa_4_87_2/B sky130_fd_sc_hd__fa_1
XFILLER_89_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_0_54_1 U$$514/X U$$647/X VGND VGND VPWR VPWR dadda_fa_1_55_8/B dadda_fa_2_54_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_2_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_57_0 dadda_fa_6_57_0/A dadda_fa_6_57_0/B dadda_fa_6_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_58_0/B dadda_fa_7_57_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_111_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4402 U$$4402/A1 U$$4388/X U$$4404/A1 U$$4508/B2 VGND VGND VPWR VPWR U$$4403/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4413 U$$4413/A U$$4413/B VGND VGND VPWR VPWR U$$4413/X sky130_fd_sc_hd__xor2_1
XU$$4424 U$$4424/A1 U$$4388/X U$$4424/B1 U$$4428/B2 VGND VGND VPWR VPWR U$$4425/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_0_60_0 U$$127/X U$$260/X U$$393/X VGND VGND VPWR VPWR dadda_fa_1_61_6/A
+ dadda_fa_1_60_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4435 U$$4435/A U$$4435/B VGND VGND VPWR VPWR U$$4435/X sky130_fd_sc_hd__xor2_1
XU$$3701 U$$3836/A VGND VGND VPWR VPWR U$$3701/Y sky130_fd_sc_hd__inv_1
XU$$4446 U$$4446/A1 U$$4388/X U$$4446/B1 U$$4506/B2 VGND VGND VPWR VPWR U$$4447/A
+ sky130_fd_sc_hd__a22o_1
XU$$3712 U$$3712/A U$$3790/B VGND VGND VPWR VPWR U$$3712/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_116_2 input147/X dadda_fa_4_116_2/B dadda_ha_3_116_0/SUM VGND VGND VPWR
+ VPWR dadda_fa_5_117_0/CIN dadda_fa_5_116_1/CIN sky130_fd_sc_hd__fa_1
XU$$4457 U$$4457/A U$$4457/B VGND VGND VPWR VPWR U$$4457/X sky130_fd_sc_hd__xor2_1
XU$$3723 U$$4132/B1 U$$3757/A2 U$$3999/A1 U$$3757/B2 VGND VGND VPWR VPWR U$$3724/A
+ sky130_fd_sc_hd__a22o_1
XU$$4468 U$$4468/A1 U$$4388/X U$$4470/A1 U$$4488/B2 VGND VGND VPWR VPWR U$$4469/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3734 U$$3734/A U$$3734/B VGND VGND VPWR VPWR U$$3734/X sky130_fd_sc_hd__xor2_1
XU$$4479 U$$4479/A U$$4479/B VGND VGND VPWR VPWR U$$4479/X sky130_fd_sc_hd__xor2_1
XU$$3745 U$$4017/B1 U$$3791/A2 U$$4432/A1 U$$3791/B2 VGND VGND VPWR VPWR U$$3746/A
+ sky130_fd_sc_hd__a22o_1
XU$$3756 U$$3756/A U$$3774/B VGND VGND VPWR VPWR U$$3756/X sky130_fd_sc_hd__xor2_1
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3767 U$$4176/B1 U$$3773/A2 U$$4043/A1 U$$3773/B2 VGND VGND VPWR VPWR U$$3768/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_109_1 dadda_fa_4_109_1/A dadda_fa_4_109_1/B dadda_fa_4_109_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_110_0/B dadda_fa_5_109_1/B sky130_fd_sc_hd__fa_1
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3778 U$$3778/A U$$3836/A VGND VGND VPWR VPWR U$$3778/X sky130_fd_sc_hd__xor2_1
XU$$3789 U$$4198/B1 U$$3791/A2 U$$4476/A1 U$$3791/B2 VGND VGND VPWR VPWR U$$3790/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_82_1 dadda_fa_2_82_1/A dadda_fa_2_82_1/B dadda_fa_2_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_0/CIN dadda_fa_3_82_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_173_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_75_0 dadda_fa_2_75_0/A dadda_fa_2_75_0/B dadda_fa_2_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_0/B dadda_fa_3_75_2/B sky130_fd_sc_hd__fa_1
XFILLER_69_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_51_7 U$$2902/X U$$3035/X U$$3168/X VGND VGND VPWR VPWR dadda_fa_2_52_2/CIN
+ dadda_fa_2_51_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3833_1825 VGND VGND VPWR VPWR U$$3833_1825/HI U$$3833/B1 sky130_fd_sc_hd__conb_1
XFILLER_110_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_97_1 dadda_fa_4_97_1/A dadda_fa_4_97_1/B dadda_fa_4_97_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_98_0/B dadda_fa_5_97_1/B sky130_fd_sc_hd__fa_1
XFILLER_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_74_0 dadda_fa_7_74_0/A dadda_fa_7_74_0/B dadda_fa_7_74_0/CIN VGND VGND
+ VPWR VPWR _371_/D _242_/D sky130_fd_sc_hd__fa_1
XFILLER_3_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1206 U$$3048/A1 VGND VGND VPWR VPWR U$$34/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1217 input68/X VGND VGND VPWR VPWR U$$4416/A1 sky130_fd_sc_hd__buf_6
XFILLER_121_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1228 U$$987/A1 VGND VGND VPWR VPWR U$$3999/B1 sky130_fd_sc_hd__buf_4
XFILLER_59_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1239 U$$828/B1 VGND VGND VPWR VPWR U$$8/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3008 U$$3008/A U$$3013/A VGND VGND VPWR VPWR U$$3008/X sky130_fd_sc_hd__xor2_1
XU$$3019 U$$3017/B U$$3014/A input39/X U$$3014/Y VGND VGND VPWR VPWR U$$3019/X sky130_fd_sc_hd__a22o_4
XFILLER_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2307 U$$2307/A U$$2329/A VGND VGND VPWR VPWR U$$2307/X sky130_fd_sc_hd__xor2_1
XU$$2318 U$$4234/B1 U$$2326/A2 U$$3964/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2319/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2329 U$$2329/A VGND VGND VPWR VPWR U$$2329/Y sky130_fd_sc_hd__inv_1
XFILLER_55_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1606 U$$1606/A U$$1608/B VGND VGND VPWR VPWR U$$1606/X sky130_fd_sc_hd__xor2_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1617 U$$521/A1 U$$1625/A2 U$$521/B1 U$$1625/B2 VGND VGND VPWR VPWR U$$1618/A sky130_fd_sc_hd__a22o_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1628 U$$1628/A U$$1630/B VGND VGND VPWR VPWR U$$1628/X sky130_fd_sc_hd__xor2_1
XU$$4465_1880 VGND VGND VPWR VPWR U$$4465_1880/HI U$$4465/B sky130_fd_sc_hd__conb_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1639 U$$4377/B1 U$$1641/A2 U$$4244/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1640/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_304_ _319_/CLK _304_/D VGND VGND VPWR VPWR _304_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_235_ _364_/CLK _235_/D VGND VGND VPWR VPWR _235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_92_0 dadda_fa_3_92_0/A dadda_fa_3_92_0/B dadda_fa_3_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_0/B dadda_fa_4_92_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1740 input104/X VGND VGND VPWR VPWR U$$783/A1 sky130_fd_sc_hd__buf_2
XFILLER_66_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1751 U$$781/A1 VGND VGND VPWR VPWR U$$3382/B1 sky130_fd_sc_hd__buf_6
Xfanout1762 U$$3243/A1 VGND VGND VPWR VPWR U$$92/A1 sky130_fd_sc_hd__buf_4
XFILLER_93_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4210 U$$4482/B1 U$$4224/A2 U$$4349/A1 U$$4224/B2 VGND VGND VPWR VPWR U$$4211/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1773 U$$3376/B1 VGND VGND VPWR VPWR U$$3239/B1 sky130_fd_sc_hd__buf_4
XFILLER_78_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_121_0 U$$3972/Y U$$4106/X U$$4239/X VGND VGND VPWR VPWR dadda_fa_5_122_1/B
+ dadda_fa_5_121_1/CIN sky130_fd_sc_hd__fa_1
XU$$4221 U$$4221/A U$$4231/B VGND VGND VPWR VPWR U$$4221/X sky130_fd_sc_hd__xor2_1
XFILLER_120_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_54_5 dadda_fa_2_54_5/A dadda_fa_2_54_5/B dadda_fa_2_54_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_2/A dadda_fa_4_54_0/A sky130_fd_sc_hd__fa_1
XFILLER_65_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4232 U$$4367/B1 U$$4236/A2 U$$4234/A1 U$$4236/B2 VGND VGND VPWR VPWR U$$4233/A
+ sky130_fd_sc_hd__a22o_1
XU$$4243 U$$4243/A U$$4247/A VGND VGND VPWR VPWR U$$4243/X sky130_fd_sc_hd__xor2_1
XU$$4254 U$$4254/A U$$4292/B VGND VGND VPWR VPWR U$$4254/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_47_4 dadda_fa_2_47_4/A dadda_fa_2_47_4/B dadda_fa_2_47_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_1/CIN dadda_fa_3_47_3/CIN sky130_fd_sc_hd__fa_1
XU$$4265 U$$4400/B1 U$$4295/A2 U$$4265/B1 U$$4295/B2 VGND VGND VPWR VPWR U$$4266/A
+ sky130_fd_sc_hd__a22o_1
XU$$3520 U$$3520/A U$$3548/B VGND VGND VPWR VPWR U$$3520/X sky130_fd_sc_hd__xor2_1
XU$$3531 U$$4214/B1 U$$3549/A2 U$$4081/A1 U$$3549/B2 VGND VGND VPWR VPWR U$$3532/A
+ sky130_fd_sc_hd__a22o_1
XU$$4276 U$$4276/A U$$4322/B VGND VGND VPWR VPWR U$$4276/X sky130_fd_sc_hd__xor2_1
XFILLER_53_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3542 U$$3542/A U$$3561/A VGND VGND VPWR VPWR U$$3542/X sky130_fd_sc_hd__xor2_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4287 U$$4287/A1 U$$4289/A2 U$$4426/A1 U$$4289/B2 VGND VGND VPWR VPWR U$$4288/A
+ sky130_fd_sc_hd__a22o_1
XU$$4298 U$$4298/A U$$4384/A VGND VGND VPWR VPWR U$$4298/X sky130_fd_sc_hd__xor2_1
XFILLER_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3553 U$$3964/A1 U$$3557/A2 U$$3966/A1 U$$3557/B2 VGND VGND VPWR VPWR U$$3554/A
+ sky130_fd_sc_hd__a22o_1
XU$$3564 U$$3699/A VGND VGND VPWR VPWR U$$3564/Y sky130_fd_sc_hd__inv_1
XFILLER_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2830 U$$3239/B1 U$$2840/A2 U$$3106/A1 U$$2840/B2 VGND VGND VPWR VPWR U$$2831/A
+ sky130_fd_sc_hd__a22o_1
XU$$3575 U$$3575/A U$$3615/B VGND VGND VPWR VPWR U$$3575/X sky130_fd_sc_hd__xor2_1
XU$$2841 U$$2841/A U$$2841/B VGND VGND VPWR VPWR U$$2841/X sky130_fd_sc_hd__xor2_1
XU$$3586 U$$4132/B1 U$$3604/A2 U$$3999/A1 U$$3604/B2 VGND VGND VPWR VPWR U$$3587/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2852 U$$4220/B1 U$$2874/A2 U$$4361/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2853/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3597 U$$3597/A U$$3601/B VGND VGND VPWR VPWR U$$3597/X sky130_fd_sc_hd__xor2_1
XU$$2863 U$$2863/A U$$2871/B VGND VGND VPWR VPWR U$$2863/X sky130_fd_sc_hd__xor2_1
XU$$2874 U$$3559/A1 U$$2874/A2 U$$2874/B1 U$$2874/B2 VGND VGND VPWR VPWR U$$2875/A
+ sky130_fd_sc_hd__a22o_1
XU$$2885 U$$3022/A1 U$$2929/A2 U$$3022/B1 U$$2929/B2 VGND VGND VPWR VPWR U$$2886/A
+ sky130_fd_sc_hd__a22o_1
XU$$2896 U$$2896/A U$$2926/B VGND VGND VPWR VPWR U$$2896/X sky130_fd_sc_hd__xor2_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_898 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$803 final_adder.U$$770/A final_adder.U$$723/X final_adder.U$$691/X
+ VGND VGND VPWR VPWR final_adder.U$$803/X sky130_fd_sc_hd__a21o_1
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$825 final_adder.U$$792/A final_adder.U$$625/X final_adder.U$$713/X
+ VGND VGND VPWR VPWR final_adder.U$$825/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$847 final_adder.U$$750/X final_adder.U$$815/X final_adder.U$$751/X
+ VGND VGND VPWR VPWR final_adder.U$$847/X sky130_fd_sc_hd__a21o_2
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$869 final_adder.U$$772/X final_adder.U$$725/X final_adder.U$$773/X
+ VGND VGND VPWR VPWR final_adder.U$$869/X sky130_fd_sc_hd__a21o_1
XU$$708 U$$708/A U$$774/B VGND VGND VPWR VPWR U$$708/X sky130_fd_sc_hd__xor2_1
XU$$719 U$$854/B1 U$$771/A2 U$$721/A1 U$$771/B2 VGND VGND VPWR VPWR U$$720/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_42_3 U$$1288/X U$$1421/X U$$1554/X VGND VGND VPWR VPWR dadda_fa_2_43_4/A
+ dadda_fa_2_42_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_12_1 U$$430/X U$$563/X U$$696/X VGND VGND VPWR VPWR dadda_fa_5_13_0/B
+ dadda_fa_5_12_1/B sky130_fd_sc_hd__fa_1
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4495_1895 VGND VGND VPWR VPWR U$$4495_1895/HI U$$4495/B sky130_fd_sc_hd__conb_1
XFILLER_106_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_109_0 U$$3150/Y U$$3284/X U$$3417/X VGND VGND VPWR VPWR dadda_fa_4_110_0/B
+ dadda_fa_4_109_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1003 U$$620/B1 VGND VGND VPWR VPWR U$$896/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1014 U$$346/A1 VGND VGND VPWR VPWR U$$72/A1 sky130_fd_sc_hd__buf_4
Xfanout1025 U$$1221/B VGND VGND VPWR VPWR U$$1175/B sky130_fd_sc_hd__buf_6
XFILLER_0_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1036 input89/X VGND VGND VPWR VPWR U$$4315/B1 sky130_fd_sc_hd__buf_6
XFILLER_66_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1047 U$$4257/B1 VGND VGND VPWR VPWR U$$3298/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_57_3 dadda_fa_3_57_3/A dadda_fa_3_57_3/B dadda_fa_3_57_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_1/B dadda_fa_4_57_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1058 U$$4450/A1 VGND VGND VPWR VPWR U$$3628/A1 sky130_fd_sc_hd__buf_6
XFILLER_102_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1069 input85/X VGND VGND VPWR VPWR U$$4446/B1 sky130_fd_sc_hd__buf_6
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2104 U$$2104/A U$$2106/B VGND VGND VPWR VPWR U$$2104/X sky130_fd_sc_hd__xor2_1
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2115 U$$745/A1 U$$2147/A2 U$$745/B1 U$$2147/B2 VGND VGND VPWR VPWR U$$2116/A sky130_fd_sc_hd__a22o_1
XU$$2126 U$$2126/A U$$2130/B VGND VGND VPWR VPWR U$$2126/X sky130_fd_sc_hd__xor2_1
XFILLER_63_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2137 U$$3642/B1 U$$2177/A2 U$$3509/A1 U$$2177/B2 VGND VGND VPWR VPWR U$$2138/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1403 U$$1403/A U$$1415/B VGND VGND VPWR VPWR U$$1403/X sky130_fd_sc_hd__xor2_1
XU$$2148 U$$2148/A U$$2148/B VGND VGND VPWR VPWR U$$2148/X sky130_fd_sc_hd__xor2_1
XFILLER_43_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2159 U$$2707/A1 U$$2177/A2 U$$2707/B1 U$$2177/B2 VGND VGND VPWR VPWR U$$2160/A
+ sky130_fd_sc_hd__a22o_1
XU$$1414 U$$316/B1 U$$1414/A2 U$$183/A1 U$$1414/B2 VGND VGND VPWR VPWR U$$1415/A sky130_fd_sc_hd__a22o_1
XU$$1425 U$$1425/A U$$1427/B VGND VGND VPWR VPWR U$$1425/X sky130_fd_sc_hd__xor2_1
XFILLER_16_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1436 U$$749/B1 U$$1452/A2 U$$616/A1 U$$1452/B2 VGND VGND VPWR VPWR U$$1437/A sky130_fd_sc_hd__a22o_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1447 U$$1447/A U$$1491/B VGND VGND VPWR VPWR U$$1447/X sky130_fd_sc_hd__xor2_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_887 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1458 U$$499/A1 U$$1460/A2 U$$90/A1 U$$1460/B2 VGND VGND VPWR VPWR U$$1459/A sky130_fd_sc_hd__a22o_1
XFILLER_163_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1469 U$$1469/A U$$1475/B VGND VGND VPWR VPWR U$$1469/X sky130_fd_sc_hd__xor2_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_218_ _218_/CLK _218_/D VGND VGND VPWR VPWR _218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_52_2 dadda_fa_2_52_2/A dadda_fa_2_52_2/B dadda_fa_2_52_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_1/A dadda_fa_3_52_3/A sky130_fd_sc_hd__fa_1
Xfanout1570 U$$3825/B1 VGND VGND VPWR VPWR U$$3964/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1581 input120/X VGND VGND VPWR VPWR U$$3580/A1 sky130_fd_sc_hd__buf_4
Xfanout1592 U$$811/A1 VGND VGND VPWR VPWR U$$672/B1 sky130_fd_sc_hd__buf_4
XU$$4040 U$$4040/A U$$4040/B VGND VGND VPWR VPWR U$$4040/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_45_1 U$$2757/X U$$2890/X U$$3023/X VGND VGND VPWR VPWR dadda_fa_3_46_0/CIN
+ dadda_fa_3_45_2/CIN sky130_fd_sc_hd__fa_1
XU$$4051 U$$4460/B1 U$$4081/A2 U$$4464/A1 U$$4081/B2 VGND VGND VPWR VPWR U$$4052/A
+ sky130_fd_sc_hd__a22o_1
XU$$4062 U$$4062/A U$$4082/B VGND VGND VPWR VPWR U$$4062/X sky130_fd_sc_hd__xor2_1
XFILLER_93_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4073 U$$4484/A1 U$$4093/A2 U$$4484/B1 U$$4093/B2 VGND VGND VPWR VPWR U$$4074/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4084 U$$4084/A U$$4098/B VGND VGND VPWR VPWR U$$4084/X sky130_fd_sc_hd__xor2_1
XU$$4095 U$$4367/B1 U$$4107/A2 U$$4234/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4096/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_22_0 dadda_fa_5_22_0/A dadda_fa_5_22_0/B dadda_fa_5_22_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_23_0/A dadda_fa_6_22_0/CIN sky130_fd_sc_hd__fa_1
XU$$3350 U$$4446/A1 U$$3416/A2 U$$4446/B1 U$$3416/B2 VGND VGND VPWR VPWR U$$3351/A
+ sky130_fd_sc_hd__a22o_1
XU$$3361 U$$3361/A U$$3373/B VGND VGND VPWR VPWR U$$3361/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_38_0 U$$1147/X U$$1280/X U$$1413/X VGND VGND VPWR VPWR dadda_fa_3_39_0/B
+ dadda_fa_3_38_2/B sky130_fd_sc_hd__fa_1
XU$$3372 U$$3509/A1 U$$3372/A2 U$$3372/B1 U$$3372/B2 VGND VGND VPWR VPWR U$$3373/A
+ sky130_fd_sc_hd__a22o_1
XU$$3383 U$$3383/A U$$3424/A VGND VGND VPWR VPWR U$$3383/X sky130_fd_sc_hd__xor2_1
XU$$3394 U$$4214/B1 U$$3416/A2 U$$4081/A1 U$$3416/B2 VGND VGND VPWR VPWR U$$3395/A
+ sky130_fd_sc_hd__a22o_1
XU$$2660 U$$2660/A U$$2662/B VGND VGND VPWR VPWR U$$2660/X sky130_fd_sc_hd__xor2_1
XU$$2671 U$$3628/B1 U$$2711/A2 U$$3630/B1 U$$2711/B2 VGND VGND VPWR VPWR U$$2672/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2682 U$$2682/A U$$2724/B VGND VGND VPWR VPWR U$$2682/X sky130_fd_sc_hd__xor2_1
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2693 U$$3239/B1 U$$2707/A2 U$$3106/A1 U$$2707/B2 VGND VGND VPWR VPWR U$$2694/A
+ sky130_fd_sc_hd__a22o_1
XU$$1970 U$$50/B1 U$$1986/A2 U$$739/A1 U$$1986/B2 VGND VGND VPWR VPWR U$$1971/A sky130_fd_sc_hd__a22o_1
XU$$1981 U$$1981/A U$$1981/B VGND VGND VPWR VPWR U$$1981/X sky130_fd_sc_hd__xor2_1
XU$$1992 U$$620/B1 U$$2006/A2 U$$898/A1 U$$2006/B2 VGND VGND VPWR VPWR U$$1993/A sky130_fd_sc_hd__a22o_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_67_2 dadda_fa_4_67_2/A dadda_fa_4_67_2/B dadda_fa_4_67_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_68_0/CIN dadda_fa_5_67_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput106 b[47] VGND VGND VPWR VPWR input106/X sky130_fd_sc_hd__buf_4
Xinput117 b[57] VGND VGND VPWR VPWR input117/X sky130_fd_sc_hd__clkbuf_1
Xinput128 b[9] VGND VGND VPWR VPWR input128/X sky130_fd_sc_hd__buf_2
Xinput139 c[109] VGND VGND VPWR VPWR input139/X sky130_fd_sc_hd__buf_2
Xfinal_adder.U$$600 final_adder.U$$608/B final_adder.U$$600/B VGND VGND VPWR VPWR
+ final_adder.U$$720/B sky130_fd_sc_hd__and2_1
XFILLER_130_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$611 final_adder.U$$610/B final_adder.U$$495/X final_adder.U$$487/X
+ VGND VGND VPWR VPWR final_adder.U$$611/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_7_37_0 dadda_fa_7_37_0/A dadda_fa_7_37_0/B dadda_fa_7_37_0/CIN VGND VGND
+ VPWR VPWR _334_/D _205_/D sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$633 final_adder.U$$632/B final_adder.U$$529/X final_adder.U$$513/X
+ VGND VGND VPWR VPWR final_adder.U$$633/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$644 final_adder.U$$660/B final_adder.U$$644/B VGND VGND VPWR VPWR
+ final_adder.U$$756/B sky130_fd_sc_hd__and2_1
XFILLER_84_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$655 final_adder.U$$654/B final_adder.U$$551/X final_adder.U$$535/X
+ VGND VGND VPWR VPWR final_adder.U$$655/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$666 final_adder.U$$682/B final_adder.U$$666/B VGND VGND VPWR VPWR
+ final_adder.U$$778/B sky130_fd_sc_hd__and2_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$505 U$$505/A1 U$$505/A2 U$$505/B1 U$$505/B2 VGND VGND VPWR VPWR U$$506/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$677 final_adder.U$$676/B final_adder.U$$573/X final_adder.U$$557/X
+ VGND VGND VPWR VPWR final_adder.U$$677/X sky130_fd_sc_hd__a21o_1
XU$$516 U$$516/A U$$522/B VGND VGND VPWR VPWR U$$516/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_40_0 U$$87/X U$$220/X U$$353/X VGND VGND VPWR VPWR dadda_fa_2_41_3/CIN
+ dadda_fa_2_40_5/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$688 final_adder.U$$704/B final_adder.U$$688/B VGND VGND VPWR VPWR
+ final_adder.U$$800/B sky130_fd_sc_hd__and2_1
XU$$527 U$$936/B1 U$$539/A2 U$$803/A1 U$$539/B2 VGND VGND VPWR VPWR U$$528/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$699 final_adder.U$$698/B final_adder.U$$595/X final_adder.U$$579/X
+ VGND VGND VPWR VPWR final_adder.U$$699/X sky130_fd_sc_hd__a21o_1
XU$$538 U$$538/A U$$548/A VGND VGND VPWR VPWR U$$538/X sky130_fd_sc_hd__xor2_1
XU$$549 U$$549/A VGND VGND VPWR VPWR U$$551/B sky130_fd_sc_hd__inv_1
XFILLER_44_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_62_1 dadda_fa_3_62_1/A dadda_fa_3_62_1/B dadda_fa_3_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_0/CIN dadda_fa_4_62_2/A sky130_fd_sc_hd__fa_1
XFILLER_79_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_55_0 dadda_fa_3_55_0/A dadda_fa_3_55_0/B dadda_fa_3_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_0/B dadda_fa_4_55_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1200 U$$2707/A1 U$$1230/A2 U$$2707/B1 U$$1230/B2 VGND VGND VPWR VPWR U$$1201/A
+ sky130_fd_sc_hd__a22o_1
XU$$1211 U$$1211/A U$$1227/B VGND VGND VPWR VPWR U$$1211/X sky130_fd_sc_hd__xor2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1222 U$$948/A1 U$$1226/A2 U$$950/A1 U$$1226/B2 VGND VGND VPWR VPWR U$$1223/A sky130_fd_sc_hd__a22o_1
XU$$1233 U$$1233/A VGND VGND VPWR VPWR U$$1233/Y sky130_fd_sc_hd__inv_1
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1244 U$$1244/A U$$1282/B VGND VGND VPWR VPWR U$$1244/X sky130_fd_sc_hd__xor2_1
XU$$1255 U$$2625/A1 U$$1295/A2 U$$983/A1 U$$1295/B2 VGND VGND VPWR VPWR U$$1256/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1266 U$$1266/A U$$1294/B VGND VGND VPWR VPWR U$$1266/X sky130_fd_sc_hd__xor2_1
XU$$1277 U$$44/A1 U$$1309/A2 U$$46/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1278/A sky130_fd_sc_hd__a22o_1
XU$$1288 U$$1288/A U$$1294/B VGND VGND VPWR VPWR U$$1288/X sky130_fd_sc_hd__xor2_1
XFILLER_148_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1299 U$$64/B1 U$$1327/A2 U$$66/B1 U$$1327/B2 VGND VGND VPWR VPWR U$$1300/A sky130_fd_sc_hd__a22o_1
XFILLER_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_112_0 dadda_fa_7_112_0/A dadda_fa_7_112_0/B dadda_fa_7_112_0/CIN VGND
+ VGND VPWR VPWR _409_/D _280_/D sky130_fd_sc_hd__fa_1
XFILLER_117_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1060 final_adder.U$$218/A final_adder.U$$831/X VGND VGND VPWR VPWR
+ output314/A sky130_fd_sc_hd__xor2_1
XFILLER_172_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1071 final_adder.U$$208/B final_adder.U$$979/X VGND VGND VPWR VPWR
+ output326/A sky130_fd_sc_hd__xor2_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1082 final_adder.U$$196/A final_adder.U$$809/X VGND VGND VPWR VPWR
+ output338/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1093 final_adder.U$$186/B final_adder.U$$957/X VGND VGND VPWR VPWR
+ output350/A sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_77_1 dadda_fa_5_77_1/A dadda_fa_5_77_1/B dadda_fa_5_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_78_0/B dadda_fa_7_77_0/A sky130_fd_sc_hd__fa_1
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout807 U$$2608/X VGND VGND VPWR VPWR U$$2711/B2 sky130_fd_sc_hd__clkbuf_4
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout818 fanout820/X VGND VGND VPWR VPWR U$$2598/B2 sky130_fd_sc_hd__buf_6
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout829 U$$2272/B2 VGND VGND VPWR VPWR U$$2254/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_8 dadda_fa_1_69_8/A dadda_fa_1_69_8/B dadda_fa_1_69_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_70_3/A dadda_fa_3_69_0/A sky130_fd_sc_hd__fa_1
XFILLER_86_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3180 U$$3180/A U$$3210/B VGND VGND VPWR VPWR U$$3180/X sky130_fd_sc_hd__xor2_1
XU$$3191 U$$4287/A1 U$$3199/A2 U$$4426/A1 U$$3199/B2 VGND VGND VPWR VPWR U$$3192/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_9_0 dadda_fa_6_9_0/A dadda_fa_6_9_0/B dadda_fa_6_9_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_10_0/B dadda_fa_7_9_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2490 U$$2762/B1 U$$2532/A2 U$$2629/A1 U$$2532/B2 VGND VGND VPWR VPWR U$$2491/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_72_0 dadda_fa_4_72_0/A dadda_fa_4_72_0/B dadda_fa_4_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_73_0/A dadda_fa_5_72_1/A sky130_fd_sc_hd__fa_1
XFILLER_116_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_88_0 dadda_fa_1_88_0/A U$$1779/X U$$1912/X VGND VGND VPWR VPWR dadda_fa_2_89_3/B
+ dadda_fa_2_88_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_107_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$430 final_adder.U$$434/B final_adder.U$$430/B VGND VGND VPWR VPWR
+ final_adder.U$$554/B sky130_fd_sc_hd__and2_1
XFILLER_29_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$441 final_adder.U$$440/B final_adder.U$$319/X final_adder.U$$315/X
+ VGND VGND VPWR VPWR final_adder.U$$441/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$452 final_adder.U$$456/B final_adder.U$$452/B VGND VGND VPWR VPWR
+ final_adder.U$$576/B sky130_fd_sc_hd__and2_1
XFILLER_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$463 final_adder.U$$462/B final_adder.U$$341/X final_adder.U$$337/X
+ VGND VGND VPWR VPWR final_adder.U$$463/X sky130_fd_sc_hd__a21o_1
XU$$302 U$$576/A1 U$$338/A2 U$$576/B1 U$$338/B2 VGND VGND VPWR VPWR U$$303/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$474 final_adder.U$$478/B final_adder.U$$474/B VGND VGND VPWR VPWR
+ final_adder.U$$598/B sky130_fd_sc_hd__and2_1
XU$$313 U$$313/A U$$313/B VGND VGND VPWR VPWR U$$313/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$485 final_adder.U$$484/B final_adder.U$$363/X final_adder.U$$359/X
+ VGND VGND VPWR VPWR final_adder.U$$485/X sky130_fd_sc_hd__a21o_1
XU$$324 U$$596/B1 U$$362/A2 U$$598/B1 U$$362/B2 VGND VGND VPWR VPWR U$$325/A sky130_fd_sc_hd__a22o_1
XFILLER_45_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$496 final_adder.U$$500/B final_adder.U$$496/B VGND VGND VPWR VPWR
+ final_adder.U$$612/A sky130_fd_sc_hd__and2_1
XFILLER_29_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$335 U$$335/A U$$353/B VGND VGND VPWR VPWR U$$335/X sky130_fd_sc_hd__xor2_1
XFILLER_45_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$346 U$$346/A1 U$$346/A2 U$$74/A1 U$$346/B2 VGND VGND VPWR VPWR U$$347/A sky130_fd_sc_hd__a22o_1
XU$$357 U$$357/A U$$363/B VGND VGND VPWR VPWR U$$357/X sky130_fd_sc_hd__xor2_1
XFILLER_26_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$368 U$$505/A1 U$$406/A2 U$$505/B1 U$$406/B2 VGND VGND VPWR VPWR U$$369/A sky130_fd_sc_hd__a22o_1
XU$$379 U$$379/A U$$387/B VGND VGND VPWR VPWR U$$379/X sky130_fd_sc_hd__xor2_1
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_87_0 dadda_fa_6_87_0/A dadda_fa_6_87_0/B dadda_fa_6_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_88_0/B dadda_fa_7_87_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_154_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3970_1827 VGND VGND VPWR VPWR U$$3970_1827/HI U$$3970/B1 sky130_fd_sc_hd__conb_1
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$880 U$$880/A1 U$$904/A2 U$$882/A1 U$$904/B2 VGND VGND VPWR VPWR U$$881/A sky130_fd_sc_hd__a22o_1
XU$$1030 U$$1030/A U$$998/B VGND VGND VPWR VPWR U$$1030/X sky130_fd_sc_hd__xor2_1
XU$$891 U$$891/A U$$895/B VGND VGND VPWR VPWR U$$891/X sky130_fd_sc_hd__xor2_1
XU$$1041 U$$82/A1 U$$981/A2 U$$82/B1 U$$981/B2 VGND VGND VPWR VPWR U$$1042/A sky130_fd_sc_hd__a22o_1
XU$$1052 U$$1052/A U$$1094/B VGND VGND VPWR VPWR U$$1052/X sky130_fd_sc_hd__xor2_1
XU$$1063 U$$926/A1 U$$963/X U$$928/A1 U$$964/X VGND VGND VPWR VPWR U$$1064/A sky130_fd_sc_hd__a22o_1
XU$$1074 U$$1074/A U$$990/B VGND VGND VPWR VPWR U$$1074/X sky130_fd_sc_hd__xor2_1
XU$$1085 U$$948/A1 U$$1087/A2 U$$950/A1 U$$1087/B2 VGND VGND VPWR VPWR U$$1086/A sky130_fd_sc_hd__a22o_1
XU$$1096 U$$962/A VGND VGND VPWR VPWR U$$1096/Y sky130_fd_sc_hd__inv_1
XFILLER_31_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_81_7 U$$4026/X U$$4159/X U$$4292/X VGND VGND VPWR VPWR dadda_fa_2_82_3/B
+ dadda_fa_3_81_0/A sky130_fd_sc_hd__fa_1
Xfanout604 U$$1726/A2 VGND VGND VPWR VPWR U$$1698/A2 sky130_fd_sc_hd__buf_2
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout615 U$$1587/A2 VGND VGND VPWR VPWR U$$1575/A2 sky130_fd_sc_hd__buf_4
XFILLER_99_985 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout626 U$$207/A2 VGND VGND VPWR VPWR U$$213/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_74_6 U$$4145/X U$$4278/X U$$4411/X VGND VGND VPWR VPWR dadda_fa_2_75_2/B
+ dadda_fa_2_74_5/B sky130_fd_sc_hd__fa_1
Xfanout637 U$$1327/A2 VGND VGND VPWR VPWR U$$1295/A2 sky130_fd_sc_hd__clkbuf_4
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout648 U$$1170/A2 VGND VGND VPWR VPWR U$$1174/A2 sky130_fd_sc_hd__buf_4
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout659 U$$964/X VGND VGND VPWR VPWR U$$1087/B2 sky130_fd_sc_hd__buf_6
XFILLER_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_67_5 input220/X dadda_fa_1_67_5/B dadda_fa_1_67_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_68_2/A dadda_fa_2_67_5/A sky130_fd_sc_hd__fa_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_957 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_62_4 U$$1727/X U$$1860/X U$$1993/X VGND VGND VPWR VPWR dadda_fa_1_63_6/CIN
+ dadda_fa_1_62_8/CIN sky130_fd_sc_hd__fa_1
XU$$3905 U$$3905/A U$$3907/B VGND VGND VPWR VPWR U$$3905/X sky130_fd_sc_hd__xor2_1
XU$$3916 U$$3916/A1 U$$3970/A2 U$$4466/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3917/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_19_2 U$$843/X U$$976/X VGND VGND VPWR VPWR dadda_fa_4_20_1/B dadda_ha_3_19_2/SUM
+ sky130_fd_sc_hd__ha_1
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$260 final_adder.U$$262/B final_adder.U$$260/B VGND VGND VPWR VPWR
+ final_adder.U$$386/B sky130_fd_sc_hd__and2_1
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3927 U$$3927/A U$$3949/B VGND VGND VPWR VPWR U$$3927/X sky130_fd_sc_hd__xor2_1
XFILLER_57_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$110 U$$521/A1 U$$120/A2 U$$521/B1 U$$120/B2 VGND VGND VPWR VPWR U$$111/A sky130_fd_sc_hd__a22o_1
XU$$3938 U$$4484/B1 U$$3960/A2 U$$4488/A1 U$$3960/B2 VGND VGND VPWR VPWR U$$3939/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$271 final_adder.U$$270/B final_adder.U$$145/X final_adder.U$$143/X
+ VGND VGND VPWR VPWR final_adder.U$$271/X sky130_fd_sc_hd__a21o_1
XFILLER_73_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3949 U$$3949/A U$$3949/B VGND VGND VPWR VPWR U$$3949/X sky130_fd_sc_hd__xor2_1
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$282 final_adder.U$$284/B final_adder.U$$282/B VGND VGND VPWR VPWR
+ final_adder.U$$408/B sky130_fd_sc_hd__and2_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_32_2 dadda_fa_3_32_2/A dadda_fa_3_32_2/B dadda_fa_3_32_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_33_1/A dadda_fa_4_32_2/B sky130_fd_sc_hd__fa_1
XU$$121 U$$121/A U$$121/B VGND VGND VPWR VPWR U$$121/X sky130_fd_sc_hd__xor2_1
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$293 final_adder.U$$292/B final_adder.U$$167/X final_adder.U$$165/X
+ VGND VGND VPWR VPWR final_adder.U$$293/X sky130_fd_sc_hd__a21o_1
XU$$132 U$$406/A1 U$$98/A2 U$$406/B1 U$$98/B2 VGND VGND VPWR VPWR U$$133/A sky130_fd_sc_hd__a22o_1
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$143 U$$143/A1 U$$179/A2 U$$965/B1 U$$179/B2 VGND VGND VPWR VPWR U$$144/A sky130_fd_sc_hd__a22o_1
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4429_1862 VGND VGND VPWR VPWR U$$4429_1862/HI U$$4429/B sky130_fd_sc_hd__conb_1
XFILLER_73_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$154 U$$154/A U$$180/B VGND VGND VPWR VPWR U$$154/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_25_1 U$$1121/X U$$1254/X U$$1387/X VGND VGND VPWR VPWR dadda_fa_4_26_0/CIN
+ dadda_fa_4_25_2/A sky130_fd_sc_hd__fa_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$165 U$$28/A1 U$$179/A2 U$$30/A1 U$$179/B2 VGND VGND VPWR VPWR U$$166/A sky130_fd_sc_hd__a22o_1
XFILLER_32_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_0__f_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _218_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$176 U$$176/A U$$210/B VGND VGND VPWR VPWR U$$176/X sky130_fd_sc_hd__xor2_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$187 U$$735/A1 U$$219/A2 U$$52/A1 U$$219/B2 VGND VGND VPWR VPWR U$$188/A sky130_fd_sc_hd__a22o_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$198 U$$198/A U$$230/B VGND VGND VPWR VPWR U$$198/X sky130_fd_sc_hd__xor2_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_18_0 U$$43/X U$$176/X U$$309/X VGND VGND VPWR VPWR dadda_fa_4_19_1/A dadda_fa_4_18_2/A
+ sky130_fd_sc_hd__fa_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_397_ _397_/CLK _397_/D VGND VGND VPWR VPWR _397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_84_5 dadda_fa_2_84_5/A dadda_fa_2_84_5/B dadda_fa_2_84_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_2/A dadda_fa_4_84_0/A sky130_fd_sc_hd__fa_2
XFILLER_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_77_4 dadda_fa_2_77_4/A dadda_fa_2_77_4/B dadda_fa_2_77_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_1/CIN dadda_fa_3_77_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_787 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2883_1812 VGND VGND VPWR VPWR U$$2883_1812/HI U$$2883/A1 sky130_fd_sc_hd__conb_1
XFILLER_64_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_100_3 U$$3665/X U$$3798/X U$$3931/X VGND VGND VPWR VPWR dadda_fa_3_101_2/B
+ dadda_fa_3_100_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_51_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_114_1 dadda_fa_5_114_1/A dadda_fa_5_114_1/B dadda_fa_5_114_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_115_0/B dadda_fa_7_114_0/A sky130_fd_sc_hd__fa_1
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_107_0 dadda_fa_5_107_0/A dadda_fa_5_107_0/B dadda_fa_5_107_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_108_0/A dadda_fa_6_107_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout401 U$$807/A2 VGND VGND VPWR VPWR U$$769/A2 sky130_fd_sc_hd__buf_4
Xfanout412 U$$638/A2 VGND VGND VPWR VPWR U$$610/A2 sky130_fd_sc_hd__buf_4
XFILLER_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_72_3 U$$3210/X U$$3343/X U$$3476/X VGND VGND VPWR VPWR dadda_fa_2_73_1/B
+ dadda_fa_2_72_4/B sky130_fd_sc_hd__fa_1
Xfanout423 U$$4309/A2 VGND VGND VPWR VPWR U$$4325/A2 sky130_fd_sc_hd__buf_6
XFILLER_132_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout434 U$$4244/A2 VGND VGND VPWR VPWR U$$4174/A2 sky130_fd_sc_hd__buf_4
Xfanout445 U$$80/A2 VGND VGND VPWR VPWR U$$48/A2 sky130_fd_sc_hd__buf_2
XFILLER_171_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout456 U$$4057/A2 VGND VGND VPWR VPWR U$$4081/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_65_2 U$$3329/X U$$3462/X U$$3595/X VGND VGND VPWR VPWR dadda_fa_2_66_1/A
+ dadda_fa_2_65_4/A sky130_fd_sc_hd__fa_1
XFILLER_48_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout467 U$$3840/X VGND VGND VPWR VPWR U$$3924/A2 sky130_fd_sc_hd__buf_6
Xfanout478 U$$3566/X VGND VGND VPWR VPWR U$$3644/A2 sky130_fd_sc_hd__buf_6
XFILLER_87_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout489 U$$3439/A2 VGND VGND VPWR VPWR U$$3549/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_42_1 dadda_fa_4_42_1/A dadda_fa_4_42_1/B dadda_fa_4_42_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_43_0/B dadda_fa_5_42_1/B sky130_fd_sc_hd__fa_1
XFILLER_111_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_58_1 U$$1985/X U$$2118/X U$$2251/X VGND VGND VPWR VPWR dadda_fa_2_59_0/CIN
+ dadda_fa_2_58_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_104_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_35_0 dadda_fa_4_35_0/A dadda_fa_4_35_0/B dadda_fa_4_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_36_0/A dadda_fa_5_35_1/A sky130_fd_sc_hd__fa_1
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_320_ _328_/CLK _320_/D VGND VGND VPWR VPWR _320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_251_ _391_/CLK _251_/D VGND VGND VPWR VPWR _251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_182_ _328_/CLK _182_/D VGND VGND VPWR VPWR _182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4459_1877 VGND VGND VPWR VPWR U$$4459_1877/HI U$$4459/B sky130_fd_sc_hd__conb_1
XFILLER_109_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_87_3 dadda_fa_3_87_3/A dadda_fa_3_87_3/B dadda_fa_3_87_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_1/B dadda_fa_4_87_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4403 U$$4403/A U$$4403/B VGND VGND VPWR VPWR U$$4403/X sky130_fd_sc_hd__xor2_1
XU$$4414 U$$4414/A1 U$$4388/X U$$4416/A1 U$$4458/B2 VGND VGND VPWR VPWR U$$4415/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_0_60_1 U$$526/X U$$659/X U$$792/X VGND VGND VPWR VPWR dadda_fa_1_61_6/B
+ dadda_fa_1_60_8/A sky130_fd_sc_hd__fa_2
XU$$4425 U$$4425/A U$$4425/B VGND VGND VPWR VPWR U$$4425/X sky130_fd_sc_hd__xor2_1
XFILLER_92_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout990 fanout993/X VGND VGND VPWR VPWR U$$215/A1 sky130_fd_sc_hd__buf_4
XU$$4436 U$$4436/A1 U$$4388/X U$$4438/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4437/A
+ sky130_fd_sc_hd__a22o_1
XU$$3702 U$$3836/A U$$3702/B VGND VGND VPWR VPWR U$$3702/X sky130_fd_sc_hd__and2_1
XU$$4447 U$$4447/A U$$4447/B VGND VGND VPWR VPWR U$$4447/X sky130_fd_sc_hd__xor2_1
XU$$3713 U$$3713/A1 U$$3739/A2 U$$3713/B1 U$$3739/B2 VGND VGND VPWR VPWR U$$3714/A
+ sky130_fd_sc_hd__a22o_1
XU$$4458 U$$4458/A1 U$$4388/X U$$4460/A1 U$$4458/B2 VGND VGND VPWR VPWR U$$4459/A
+ sky130_fd_sc_hd__a22o_1
XU$$3724 U$$3724/A U$$3734/B VGND VGND VPWR VPWR U$$3724/X sky130_fd_sc_hd__xor2_1
XU$$4469 U$$4469/A U$$4469/B VGND VGND VPWR VPWR U$$4469/X sky130_fd_sc_hd__xor2_1
XU$$3735 U$$3870/B1 U$$3739/A2 U$$4420/B1 U$$3739/B2 VGND VGND VPWR VPWR U$$3736/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_161_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3746 U$$3746/A U$$3790/B VGND VGND VPWR VPWR U$$3746/X sky130_fd_sc_hd__xor2_1
XU$$3757 U$$4442/A1 U$$3757/A2 U$$4442/B1 U$$3757/B2 VGND VGND VPWR VPWR U$$3758/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3768 U$$3768/A U$$3774/B VGND VGND VPWR VPWR U$$3768/X sky130_fd_sc_hd__xor2_1
XFILLER_18_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_109_2 dadda_fa_4_109_2/A dadda_fa_4_109_2/B dadda_fa_4_109_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_110_0/CIN dadda_fa_5_109_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3779 U$$3916/A1 U$$3829/A2 U$$4466/A1 U$$3829/B2 VGND VGND VPWR VPWR U$$3780/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_82_2 dadda_fa_2_82_2/A dadda_fa_2_82_2/B dadda_fa_2_82_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_1/A dadda_fa_3_82_3/A sky130_fd_sc_hd__fa_1
XFILLER_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_75_1 dadda_fa_2_75_1/A dadda_fa_2_75_1/B dadda_fa_2_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_0/CIN dadda_fa_3_75_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_52_0 dadda_fa_5_52_0/A dadda_fa_5_52_0/B dadda_fa_5_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_53_0/A dadda_fa_6_52_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_2_68_0 dadda_fa_2_68_0/A dadda_fa_2_68_0/B dadda_fa_2_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_0/B dadda_fa_3_68_2/B sky130_fd_sc_hd__fa_1
XFILLER_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_919 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_97_2 dadda_fa_4_97_2/A dadda_fa_4_97_2/B dadda_fa_4_97_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_98_0/CIN dadda_fa_5_97_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_166_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_67_0 dadda_fa_7_67_0/A dadda_fa_7_67_0/B dadda_fa_7_67_0/CIN VGND VGND
+ VPWR VPWR _364_/D _235_/D sky130_fd_sc_hd__fa_1
XFILLER_8_1011 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1207 U$$3048/A1 VGND VGND VPWR VPWR U$$32/B1 sky130_fd_sc_hd__buf_4
Xfanout1218 U$$2631/B1 VGND VGND VPWR VPWR U$$989/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_70_0 U$$2275/X U$$2408/X U$$2541/X VGND VGND VPWR VPWR dadda_fa_2_71_0/B
+ dadda_fa_2_70_3/B sky130_fd_sc_hd__fa_1
Xfanout1229 input66/X VGND VGND VPWR VPWR U$$987/A1 sky130_fd_sc_hd__buf_4
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3009 U$$3418/B1 U$$3011/A2 U$$3285/A1 U$$3011/B2 VGND VGND VPWR VPWR U$$3010/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2308 U$$2443/B1 U$$2310/A2 U$$2310/A1 U$$2310/B2 VGND VGND VPWR VPWR U$$2309/A
+ sky130_fd_sc_hd__a22o_1
XU$$2319 U$$2319/A U$$2328/A VGND VGND VPWR VPWR U$$2319/X sky130_fd_sc_hd__xor2_1
XFILLER_28_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1607 U$$98/B1 U$$1641/A2 U$$924/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1608/A sky130_fd_sc_hd__a22o_1
XFILLER_54_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1618 U$$1618/A U$$1618/B VGND VGND VPWR VPWR U$$1618/X sky130_fd_sc_hd__xor2_1
XFILLER_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1629 U$$2175/B1 U$$1641/A2 U$$2042/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1630/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_303_ _319_/CLK _303_/D VGND VGND VPWR VPWR _303_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_234_ _364_/CLK _234_/D VGND VGND VPWR VPWR _234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_92_1 dadda_fa_3_92_1/A dadda_fa_3_92_1/B dadda_fa_3_92_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_0/CIN dadda_fa_4_92_2/A sky130_fd_sc_hd__fa_1
XFILLER_109_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_85_0 dadda_fa_3_85_0/A dadda_fa_3_85_0/B dadda_fa_3_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_0/B dadda_fa_4_85_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_123_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1730 input105/X VGND VGND VPWR VPWR U$$920/B1 sky130_fd_sc_hd__buf_6
Xfanout1741 U$$3249/A1 VGND VGND VPWR VPWR U$$4345/A1 sky130_fd_sc_hd__buf_4
Xfanout1752 input103/X VGND VGND VPWR VPWR U$$781/A1 sky130_fd_sc_hd__buf_4
XU$$4200 U$$4474/A1 U$$4226/A2 U$$4474/B1 U$$4226/B2 VGND VGND VPWR VPWR U$$4201/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_172_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1763 U$$3243/A1 VGND VGND VPWR VPWR U$$503/A1 sky130_fd_sc_hd__buf_4
XU$$4211 U$$4211/A U$$4215/B VGND VGND VPWR VPWR U$$4211/X sky130_fd_sc_hd__xor2_1
Xfanout1774 input100/X VGND VGND VPWR VPWR U$$3376/B1 sky130_fd_sc_hd__buf_6
XU$$4222 U$$4359/A1 U$$4226/A2 U$$4359/B1 U$$4226/B2 VGND VGND VPWR VPWR U$$4223/A
+ sky130_fd_sc_hd__a22o_1
XU$$4233 U$$4233/A U$$4241/B VGND VGND VPWR VPWR U$$4233/X sky130_fd_sc_hd__xor2_1
XFILLER_120_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4244 U$$4244/A1 U$$4244/A2 U$$4244/B1 U$$4244/B2 VGND VGND VPWR VPWR U$$4245/A
+ sky130_fd_sc_hd__a22o_1
XU$$3510 U$$3510/A U$$3562/A VGND VGND VPWR VPWR U$$3510/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_47_5 dadda_fa_2_47_5/A dadda_fa_2_47_5/B dadda_fa_2_47_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_2/A dadda_fa_4_47_0/A sky130_fd_sc_hd__fa_1
XU$$4255 U$$4392/A1 U$$4295/A2 U$$4257/A1 U$$4295/B2 VGND VGND VPWR VPWR U$$4256/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_114_0 U$$4092/X U$$4225/X U$$4358/X VGND VGND VPWR VPWR dadda_fa_5_115_0/A
+ dadda_fa_5_114_1/A sky130_fd_sc_hd__fa_1
XU$$4266 U$$4266/A U$$4292/B VGND VGND VPWR VPWR U$$4266/X sky130_fd_sc_hd__xor2_1
XU$$3521 U$$918/A1 U$$3523/A2 U$$920/A1 U$$3523/B2 VGND VGND VPWR VPWR U$$3522/A sky130_fd_sc_hd__a22o_1
XU$$3532 U$$3532/A U$$3548/B VGND VGND VPWR VPWR U$$3532/X sky130_fd_sc_hd__xor2_1
XU$$4277 U$$4414/A1 U$$4325/A2 U$$4416/A1 U$$4325/B2 VGND VGND VPWR VPWR U$$4278/A
+ sky130_fd_sc_hd__a22o_1
XU$$4288 U$$4288/A U$$4292/B VGND VGND VPWR VPWR U$$4288/X sky130_fd_sc_hd__xor2_1
XU$$3543 U$$4226/B1 U$$3559/A2 U$$4093/A1 U$$3559/B2 VGND VGND VPWR VPWR U$$3544/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3554 U$$3554/A U$$3558/B VGND VGND VPWR VPWR U$$3554/X sky130_fd_sc_hd__xor2_1
XU$$4299 U$$4436/A1 U$$4381/A2 U$$4438/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4300/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2820 U$$3916/A1 U$$2872/A2 U$$4464/B1 U$$2872/B2 VGND VGND VPWR VPWR U$$2821/A
+ sky130_fd_sc_hd__a22o_1
XU$$3565 U$$3699/A U$$3565/B VGND VGND VPWR VPWR U$$3565/X sky130_fd_sc_hd__and2_1
XU$$2831 U$$2831/A U$$2841/B VGND VGND VPWR VPWR U$$2831/X sky130_fd_sc_hd__xor2_1
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3576 U$$3713/A1 U$$3656/A2 U$$3713/B1 U$$3656/B2 VGND VGND VPWR VPWR U$$3577/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3587 U$$3587/A U$$3601/B VGND VGND VPWR VPWR U$$3587/X sky130_fd_sc_hd__xor2_1
XU$$2842 U$$922/B1 U$$2844/A2 U$$2979/B1 U$$2844/B2 VGND VGND VPWR VPWR U$$2843/A
+ sky130_fd_sc_hd__a22o_1
XU$$3598 U$$3870/B1 U$$3604/A2 U$$4420/B1 U$$3604/B2 VGND VGND VPWR VPWR U$$3599/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2853 U$$2853/A U$$2876/A VGND VGND VPWR VPWR U$$2853/X sky130_fd_sc_hd__xor2_1
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2864 U$$3684/B1 U$$2874/A2 U$$3551/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2865/A
+ sky130_fd_sc_hd__a22o_1
XU$$2875 U$$2875/A U$$2876/A VGND VGND VPWR VPWR U$$2875/X sky130_fd_sc_hd__xor2_1
XU$$2886 U$$2886/A U$$2926/B VGND VGND VPWR VPWR U$$2886/X sky130_fd_sc_hd__xor2_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2897 U$$2897/A1 U$$2937/A2 U$$2897/B1 U$$2937/B2 VGND VGND VPWR VPWR U$$2898/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$815 final_adder.U$$782/A final_adder.U$$735/X final_adder.U$$703/X
+ VGND VGND VPWR VPWR final_adder.U$$815/X sky130_fd_sc_hd__a21o_1
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$837 final_adder.U$$740/X final_adder.U$$805/X final_adder.U$$741/X
+ VGND VGND VPWR VPWR final_adder.U$$837/X sky130_fd_sc_hd__a21o_4
Xfinal_adder.U$$859 final_adder.U$$762/X final_adder.U$$827/X final_adder.U$$763/X
+ VGND VGND VPWR VPWR final_adder.U$$859/X sky130_fd_sc_hd__a21o_1
XU$$709 U$$709/A1 U$$743/A2 U$$709/B1 U$$743/B2 VGND VGND VPWR VPWR U$$710/A sky130_fd_sc_hd__a22o_1
XFILLER_83_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_109_1 U$$3550/X U$$3683/X U$$3816/X VGND VGND VPWR VPWR dadda_fa_4_110_0/CIN
+ dadda_fa_4_109_2/A sky130_fd_sc_hd__fa_1
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1004 fanout1011/X VGND VGND VPWR VPWR U$$620/B1 sky130_fd_sc_hd__buf_4
XFILLER_117_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1015 U$$4182/A1 VGND VGND VPWR VPWR U$$346/A1 sky130_fd_sc_hd__buf_4
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1026 U$$1221/B VGND VGND VPWR VPWR U$$1171/B sky130_fd_sc_hd__buf_6
Xfanout1037 U$$68/A1 VGND VGND VPWR VPWR U$$66/B1 sky130_fd_sc_hd__buf_4
Xfanout1048 U$$4396/A1 VGND VGND VPWR VPWR U$$4257/B1 sky130_fd_sc_hd__buf_4
XFILLER_102_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1059 U$$4450/A1 VGND VGND VPWR VPWR U$$4176/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2105 U$$872/A1 U$$2147/A2 U$$874/A1 U$$2147/B2 VGND VGND VPWR VPWR U$$2106/A sky130_fd_sc_hd__a22o_1
XFILLER_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2116 U$$2116/A U$$2148/B VGND VGND VPWR VPWR U$$2116/X sky130_fd_sc_hd__xor2_1
XU$$2127 U$$70/B1 U$$2139/A2 U$$620/B1 U$$2139/B2 VGND VGND VPWR VPWR U$$2128/A sky130_fd_sc_hd__a22o_1
XU$$2138 U$$2138/A U$$2168/B VGND VGND VPWR VPWR U$$2138/X sky130_fd_sc_hd__xor2_1
XU$$1404 U$$32/B1 U$$1414/A2 U$$447/A1 U$$1414/B2 VGND VGND VPWR VPWR U$$1405/A sky130_fd_sc_hd__a22o_1
XU$$2149 U$$916/A1 U$$2189/A2 U$$918/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2150/A sky130_fd_sc_hd__a22o_1
XU$$1415 U$$1415/A U$$1415/B VGND VGND VPWR VPWR U$$1415/X sky130_fd_sc_hd__xor2_1
XFILLER_27_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1426 U$$465/B1 U$$1426/A2 U$$58/A1 U$$1426/B2 VGND VGND VPWR VPWR U$$1427/A sky130_fd_sc_hd__a22o_1
XU$$1437 U$$1437/A U$$1449/B VGND VGND VPWR VPWR U$$1437/X sky130_fd_sc_hd__xor2_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1448 U$$78/A1 U$$1480/A2 U$$80/A1 U$$1480/B2 VGND VGND VPWR VPWR U$$1449/A sky130_fd_sc_hd__a22o_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1459 U$$1459/A U$$1461/B VGND VGND VPWR VPWR U$$1459/X sky130_fd_sc_hd__xor2_1
XFILLER_16_899 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_217_ _345_/CLK _217_/D VGND VGND VPWR VPWR _217_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_11_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1560 U$$3692/A1 VGND VGND VPWR VPWR U$$3966/A1 sky130_fd_sc_hd__buf_2
Xdadda_fa_2_52_3 dadda_fa_2_52_3/A dadda_fa_2_52_3/B dadda_fa_2_52_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_1/B dadda_fa_3_52_3/B sky130_fd_sc_hd__fa_1
Xfanout1571 U$$3825/B1 VGND VGND VPWR VPWR U$$3416/A1 sky130_fd_sc_hd__buf_4
XU$$4030 U$$4030/A U$$4040/B VGND VGND VPWR VPWR U$$4030/X sky130_fd_sc_hd__xor2_1
Xfanout1582 U$$127/B VGND VGND VPWR VPWR U$$97/B sky130_fd_sc_hd__buf_6
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4041 U$$4176/B1 U$$4043/A2 U$$4043/A1 U$$4043/B2 VGND VGND VPWR VPWR U$$4042/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1593 U$$811/A1 VGND VGND VPWR VPWR U$$2179/B1 sky130_fd_sc_hd__buf_4
XU$$4052 U$$4052/A U$$4082/B VGND VGND VPWR VPWR U$$4052/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_45_2 input196/X dadda_fa_2_45_2/B dadda_fa_2_45_2/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_46_1/A dadda_fa_3_45_3/A sky130_fd_sc_hd__fa_1
XU$$4063 U$$4198/B1 U$$4081/A2 U$$4476/A1 U$$4081/B2 VGND VGND VPWR VPWR U$$4064/A
+ sky130_fd_sc_hd__a22o_1
XU$$4074 U$$4074/A U$$4094/B VGND VGND VPWR VPWR U$$4074/X sky130_fd_sc_hd__xor2_1
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3340 U$$874/A1 U$$3340/A2 U$$876/A1 U$$3340/B2 VGND VGND VPWR VPWR U$$3341/A sky130_fd_sc_hd__a22o_1
XFILLER_93_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4085 U$$4220/B1 U$$4105/A2 U$$4361/A1 U$$4105/B2 VGND VGND VPWR VPWR U$$4086/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_22_1 dadda_fa_5_22_1/A dadda_fa_5_22_1/B dadda_fa_5_22_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_23_0/B dadda_fa_7_22_0/A sky130_fd_sc_hd__fa_1
XFILLER_53_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4096 U$$4096/A U$$4098/B VGND VGND VPWR VPWR U$$4096/X sky130_fd_sc_hd__xor2_1
XU$$3351 U$$3351/A U$$3417/B VGND VGND VPWR VPWR U$$3351/X sky130_fd_sc_hd__xor2_1
XFILLER_25_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3362 U$$3499/A1 U$$3372/A2 U$$3636/B1 U$$3372/B2 VGND VGND VPWR VPWR U$$3363/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_38_1 U$$1546/X U$$1679/X U$$1812/X VGND VGND VPWR VPWR dadda_fa_3_39_0/CIN
+ dadda_fa_3_38_2/CIN sky130_fd_sc_hd__fa_1
XU$$3373 U$$3373/A U$$3373/B VGND VGND VPWR VPWR U$$3373/X sky130_fd_sc_hd__xor2_1
XFILLER_65_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3384 U$$4478/B1 U$$3422/A2 U$$4345/A1 U$$3422/B2 VGND VGND VPWR VPWR U$$3385/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_45_clk _218_/CLK VGND VGND VPWR VPWR _343_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_5_15_0 dadda_fa_5_15_0/A dadda_fa_5_15_0/B dadda_fa_5_15_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_16_0/A dadda_fa_6_15_0/CIN sky130_fd_sc_hd__fa_2
XU$$3395 U$$3395/A U$$3417/B VGND VGND VPWR VPWR U$$3395/X sky130_fd_sc_hd__xor2_1
XU$$2650 U$$2650/A U$$2678/B VGND VGND VPWR VPWR U$$2650/X sky130_fd_sc_hd__xor2_1
XU$$2661 U$$3072/A1 U$$2667/A2 U$$3072/B1 U$$2667/B2 VGND VGND VPWR VPWR U$$2662/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2672 U$$2672/A U$$2740/A VGND VGND VPWR VPWR U$$2672/X sky130_fd_sc_hd__xor2_1
XFILLER_33_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2683 U$$3916/A1 U$$2733/A2 U$$4464/B1 U$$2733/B2 VGND VGND VPWR VPWR U$$2684/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2694 U$$2694/A U$$2708/B VGND VGND VPWR VPWR U$$2694/X sky130_fd_sc_hd__xor2_1
XFILLER_90_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1960 U$$3056/A1 U$$1964/A2 U$$3056/B1 U$$1964/B2 VGND VGND VPWR VPWR U$$1961/A
+ sky130_fd_sc_hd__a22o_1
XU$$1971 U$$1971/A U$$1971/B VGND VGND VPWR VPWR U$$1971/X sky130_fd_sc_hd__xor2_1
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1982 U$$612/A1 U$$2014/A2 U$$612/B1 U$$2014/B2 VGND VGND VPWR VPWR U$$1983/A sky130_fd_sc_hd__a22o_1
XU$$1993 U$$1993/A U$$2007/B VGND VGND VPWR VPWR U$$1993/X sky130_fd_sc_hd__xor2_1
XFILLER_21_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_41_3 U$$1286/X U$$1419/X VGND VGND VPWR VPWR dadda_fa_2_42_4/B dadda_fa_3_41_0/A
+ sky130_fd_sc_hd__ha_1
Xinput107 b[48] VGND VGND VPWR VPWR input107/X sky130_fd_sc_hd__clkbuf_1
Xinput118 b[58] VGND VGND VPWR VPWR input118/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput129 c[0] VGND VGND VPWR VPWR _296_/D sky130_fd_sc_hd__clkbuf_4
Xfinal_adder.U$$601 final_adder.U$$600/B final_adder.U$$485/X final_adder.U$$477/X
+ VGND VGND VPWR VPWR final_adder.U$$601/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$612 final_adder.U$$612/A final_adder.U$$612/B VGND VGND VPWR VPWR
+ final_adder.U$$716/A sky130_fd_sc_hd__and2_1
XFILLER_130_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$623 final_adder.U$$614/A final_adder.U$$381/X final_adder.U$$499/X
+ VGND VGND VPWR VPWR final_adder.U$$623/X sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$634 final_adder.U$$650/B final_adder.U$$634/B VGND VGND VPWR VPWR
+ final_adder.U$$746/B sky130_fd_sc_hd__and2_1
XFILLER_111_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_4_11_1 U$$428/X U$$561/X VGND VGND VPWR VPWR dadda_fa_5_12_0/CIN dadda_ha_4_11_1/SUM
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$645 final_adder.U$$644/B final_adder.U$$541/X final_adder.U$$525/X
+ VGND VGND VPWR VPWR final_adder.U$$645/X sky130_fd_sc_hd__a21o_1
XFILLER_29_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$656 final_adder.U$$672/B final_adder.U$$656/B VGND VGND VPWR VPWR
+ final_adder.U$$768/B sky130_fd_sc_hd__and2_1
XFILLER_84_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$667 final_adder.U$$666/B final_adder.U$$563/X final_adder.U$$547/X
+ VGND VGND VPWR VPWR final_adder.U$$667/X sky130_fd_sc_hd__a21o_1
XU$$506 U$$506/A U$$506/B VGND VGND VPWR VPWR U$$506/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$678 final_adder.U$$694/B final_adder.U$$678/B VGND VGND VPWR VPWR
+ final_adder.U$$790/B sky130_fd_sc_hd__and2_1
XU$$517 U$$517/A1 U$$545/A2 U$$517/B1 U$$545/B2 VGND VGND VPWR VPWR U$$518/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$689 final_adder.U$$688/B final_adder.U$$585/X final_adder.U$$569/X
+ VGND VGND VPWR VPWR final_adder.U$$689/X sky130_fd_sc_hd__a21o_1
XU$$528 U$$528/A U$$536/B VGND VGND VPWR VPWR U$$528/X sky130_fd_sc_hd__xor2_1
XFILLER_44_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_40_1 U$$486/X U$$619/X U$$752/X VGND VGND VPWR VPWR dadda_fa_2_41_4/A
+ dadda_fa_2_40_5/B sky130_fd_sc_hd__fa_1
XFILLER_16_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$539 U$$539/A1 U$$539/A2 U$$539/B1 U$$539/B2 VGND VGND VPWR VPWR U$$540/A sky130_fd_sc_hd__a22o_1
XFILLER_44_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_36_clk _388_/CLK VGND VGND VPWR VPWR _380_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_62_2 dadda_fa_3_62_2/A dadda_fa_3_62_2/B dadda_fa_3_62_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_1/A dadda_fa_4_62_2/B sky130_fd_sc_hd__fa_1
XFILLER_79_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_55_1 dadda_fa_3_55_1/A dadda_fa_3_55_1/B dadda_fa_3_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_0/CIN dadda_fa_4_55_2/A sky130_fd_sc_hd__fa_1
XFILLER_130_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_32_0 dadda_fa_6_32_0/A dadda_fa_6_32_0/B dadda_fa_6_32_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_33_0/B dadda_fa_7_32_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_48_0 dadda_fa_3_48_0/A dadda_fa_3_48_0/B dadda_fa_3_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_0/B dadda_fa_4_48_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_clk _388_/CLK VGND VGND VPWR VPWR _422_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1201 U$$1201/A U$$1233/A VGND VGND VPWR VPWR U$$1201/X sky130_fd_sc_hd__xor2_1
XU$$1212 U$$253/A1 U$$1226/A2 U$$253/B1 U$$1226/B2 VGND VGND VPWR VPWR U$$1213/A sky130_fd_sc_hd__a22o_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1223 U$$1223/A U$$1227/B VGND VGND VPWR VPWR U$$1223/X sky130_fd_sc_hd__xor2_1
XU$$1234 input10/X VGND VGND VPWR VPWR U$$1236/B sky130_fd_sc_hd__inv_1
XFILLER_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1245 U$$697/A1 U$$1309/A2 U$$697/B1 U$$1309/B2 VGND VGND VPWR VPWR U$$1246/A sky130_fd_sc_hd__a22o_1
XU$$1256 U$$1256/A U$$1294/B VGND VGND VPWR VPWR U$$1256/X sky130_fd_sc_hd__xor2_1
XU$$1267 U$$854/B1 U$$1311/A2 U$$3322/B1 U$$1311/B2 VGND VGND VPWR VPWR U$$1268/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1278 U$$1278/A U$$1278/B VGND VGND VPWR VPWR U$$1278/X sky130_fd_sc_hd__xor2_1
XU$$1289 U$$465/B1 U$$1295/A2 U$$58/A1 U$$1295/B2 VGND VGND VPWR VPWR U$$1290/A sky130_fd_sc_hd__a22o_1
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_105_0 dadda_fa_7_105_0/A dadda_fa_7_105_0/B dadda_fa_7_105_0/CIN VGND
+ VGND VPWR VPWR _402_/D _273_/D sky130_fd_sc_hd__fa_1
XFILLER_157_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1050 final_adder.U$$228/A final_adder.U$$729/X VGND VGND VPWR VPWR
+ output303/A sky130_fd_sc_hd__xor2_1
XFILLER_8_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1061 final_adder.U$$218/B final_adder.U$$989/X VGND VGND VPWR VPWR
+ output315/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1072 final_adder.U$$206/A final_adder.U$$819/X VGND VGND VPWR VPWR
+ output327/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1083 final_adder.U$$196/B final_adder.U$$967/X VGND VGND VPWR VPWR
+ output339/A sky130_fd_sc_hd__xor2_1
XFILLER_172_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1094 final_adder.U$$184/A final_adder.U$$893/X VGND VGND VPWR VPWR
+ output352/A sky130_fd_sc_hd__xor2_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout808 U$$2679/B2 VGND VGND VPWR VPWR U$$2681/B2 sky130_fd_sc_hd__buf_6
Xfanout819 fanout820/X VGND VGND VPWR VPWR U$$2600/B2 sky130_fd_sc_hd__clkbuf_4
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_50_0 U$$3474/B input202/X dadda_fa_2_50_0/CIN VGND VGND VPWR VPWR dadda_fa_3_51_0/B
+ dadda_fa_3_50_2/B sky130_fd_sc_hd__fa_1
Xfanout1390 fanout1391/X VGND VGND VPWR VPWR U$$2873/B sky130_fd_sc_hd__buf_6
XFILLER_54_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_clk _370_/CLK VGND VGND VPWR VPWR _420_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$3170 U$$3170/A U$$3210/B VGND VGND VPWR VPWR U$$3170/X sky130_fd_sc_hd__xor2_1
XU$$3181 U$$3181/A1 U$$3255/A2 U$$3181/B1 U$$3255/B2 VGND VGND VPWR VPWR U$$3182/A
+ sky130_fd_sc_hd__a22o_1
XU$$3192 U$$3192/A U$$3196/B VGND VGND VPWR VPWR U$$3192/X sky130_fd_sc_hd__xor2_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2480 U$$2480/A1 U$$2540/A2 U$$3850/B1 U$$2540/B2 VGND VGND VPWR VPWR U$$2481/A
+ sky130_fd_sc_hd__a22o_1
XU$$2491 U$$2491/A U$$2529/B VGND VGND VPWR VPWR U$$2491/X sky130_fd_sc_hd__xor2_1
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1790 U$$1790/A U$$1828/B VGND VGND VPWR VPWR U$$1790/X sky130_fd_sc_hd__xor2_1
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_72_1 dadda_fa_4_72_1/A dadda_fa_4_72_1/B dadda_fa_4_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_73_0/B dadda_fa_5_72_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_88_1 U$$2045/X U$$2178/X U$$2311/X VGND VGND VPWR VPWR dadda_fa_2_89_3/CIN
+ dadda_fa_2_88_5/A sky130_fd_sc_hd__fa_1
XFILLER_107_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_65_0 dadda_fa_4_65_0/A dadda_fa_4_65_0/B dadda_fa_4_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_66_0/A dadda_fa_5_65_1/A sky130_fd_sc_hd__fa_1
XFILLER_1_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$420 final_adder.U$$424/B final_adder.U$$420/B VGND VGND VPWR VPWR
+ final_adder.U$$544/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$431 final_adder.U$$430/B final_adder.U$$309/X final_adder.U$$305/X
+ VGND VGND VPWR VPWR final_adder.U$$431/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$442 final_adder.U$$446/B final_adder.U$$442/B VGND VGND VPWR VPWR
+ final_adder.U$$566/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$453 final_adder.U$$452/B final_adder.U$$331/X final_adder.U$$327/X
+ VGND VGND VPWR VPWR final_adder.U$$453/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$464 final_adder.U$$468/B final_adder.U$$464/B VGND VGND VPWR VPWR
+ final_adder.U$$588/B sky130_fd_sc_hd__and2_1
XU$$303 U$$303/A U$$339/B VGND VGND VPWR VPWR U$$303/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$475 final_adder.U$$474/B final_adder.U$$353/X final_adder.U$$349/X
+ VGND VGND VPWR VPWR final_adder.U$$475/X sky130_fd_sc_hd__a21o_1
XFILLER_83_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$314 U$$314/A1 U$$340/A2 U$$42/A1 U$$340/B2 VGND VGND VPWR VPWR U$$315/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$486 final_adder.U$$490/B final_adder.U$$486/B VGND VGND VPWR VPWR
+ final_adder.U$$610/B sky130_fd_sc_hd__and2_1
XU$$325 U$$325/A U$$363/B VGND VGND VPWR VPWR U$$325/X sky130_fd_sc_hd__xor2_1
XFILLER_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$497 final_adder.U$$496/B final_adder.U$$375/X final_adder.U$$371/X
+ VGND VGND VPWR VPWR final_adder.U$$497/X sky130_fd_sc_hd__a21o_1
XFILLER_44_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$336 U$$884/A1 U$$352/A2 U$$884/B1 U$$352/B2 VGND VGND VPWR VPWR U$$337/A sky130_fd_sc_hd__a22o_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$347 U$$347/A U$$347/B VGND VGND VPWR VPWR U$$347/X sky130_fd_sc_hd__xor2_1
XU$$358 U$$632/A1 U$$362/A2 U$$632/B1 U$$362/B2 VGND VGND VPWR VPWR U$$359/A sky130_fd_sc_hd__a22o_1
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$369 U$$369/A U$$407/B VGND VGND VPWR VPWR U$$369/X sky130_fd_sc_hd__xor2_1
XFILLER_26_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$870 U$$870/A1 U$$876/A2 U$$872/A1 U$$876/B2 VGND VGND VPWR VPWR U$$871/A sky130_fd_sc_hd__a22o_1
XU$$1020 U$$1020/A U$$1062/B VGND VGND VPWR VPWR U$$1020/X sky130_fd_sc_hd__xor2_1
XU$$881 U$$881/A U$$907/B VGND VGND VPWR VPWR U$$881/X sky130_fd_sc_hd__xor2_1
XU$$892 U$$892/A1 U$$898/A2 U$$894/A1 U$$898/B2 VGND VGND VPWR VPWR U$$893/A sky130_fd_sc_hd__a22o_1
XU$$1031 U$$894/A1 U$$999/A2 U$$896/A1 U$$999/B2 VGND VGND VPWR VPWR U$$1032/A sky130_fd_sc_hd__a22o_1
XU$$1042 U$$1042/A U$$1046/B VGND VGND VPWR VPWR U$$1042/X sky130_fd_sc_hd__xor2_1
XU$$1053 U$$916/A1 U$$1093/A2 U$$918/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1054/A sky130_fd_sc_hd__a22o_1
XU$$1064 U$$1064/A U$$962/A VGND VGND VPWR VPWR U$$1064/X sky130_fd_sc_hd__xor2_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1075 U$$936/B1 U$$1075/A2 U$$803/A1 U$$1075/B2 VGND VGND VPWR VPWR U$$1076/A sky130_fd_sc_hd__a22o_1
XU$$1086 U$$1086/A U$$1088/B VGND VGND VPWR VPWR U$$1086/X sky130_fd_sc_hd__xor2_1
XU$$1097 input8/X VGND VGND VPWR VPWR U$$1099/B sky130_fd_sc_hd__inv_1
XFILLER_31_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_82_0 dadda_fa_5_82_0/A dadda_fa_5_82_0/B dadda_fa_5_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_83_0/A dadda_fa_6_82_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_98_0 dadda_fa_2_98_0/A U$$2464/X U$$2597/X VGND VGND VPWR VPWR dadda_fa_3_99_0/CIN
+ dadda_fa_3_98_2/B sky130_fd_sc_hd__fa_1
XFILLER_144_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_clk _201_/CLK VGND VGND VPWR VPWR _353_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout605 U$$1760/A2 VGND VGND VPWR VPWR U$$1726/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout616 U$$1621/A2 VGND VGND VPWR VPWR U$$1587/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout627 U$$253/A2 VGND VGND VPWR VPWR U$$207/A2 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_1_74_7 input228/X dadda_fa_1_74_7/B dadda_fa_1_74_7/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_75_2/CIN dadda_fa_2_74_5/CIN sky130_fd_sc_hd__fa_1
Xfanout638 U$$1361/A2 VGND VGND VPWR VPWR U$$1327/A2 sky130_fd_sc_hd__buf_4
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout649 U$$1218/A2 VGND VGND VPWR VPWR U$$1170/A2 sky130_fd_sc_hd__buf_4
XFILLER_100_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_6 dadda_fa_1_67_6/A dadda_fa_1_67_6/B dadda_fa_1_67_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_68_2/B dadda_fa_2_67_5/B sky130_fd_sc_hd__fa_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_1_94_1 U$$2456/X U$$2589/X VGND VGND VPWR VPWR dadda_fa_2_95_5/CIN dadda_fa_3_94_0/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_7_97_0 dadda_fa_7_97_0/A dadda_fa_7_97_0/B dadda_fa_7_97_0/CIN VGND VGND
+ VPWR VPWR _394_/D _265_/D sky130_fd_sc_hd__fa_1
XFILLER_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_112_0 dadda_fa_6_112_0/A dadda_fa_6_112_0/B dadda_fa_6_112_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_113_0/B dadda_fa_7_112_0/CIN sky130_fd_sc_hd__fa_1
XU$$3906 U$$4043/A1 U$$3906/A2 U$$4043/B1 U$$3906/B2 VGND VGND VPWR VPWR U$$3907/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3917 U$$3917/A U$$3965/B VGND VGND VPWR VPWR U$$3917/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$250 final_adder.U$$4/SUM final_adder.U$$5/SUM VGND VGND VPWR VPWR
+ final_adder.U$$378/B sky130_fd_sc_hd__and2_1
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3928 U$$4474/B1 U$$3948/A2 U$$4341/A1 U$$3948/B2 VGND VGND VPWR VPWR U$$3929/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$261 final_adder.U$$260/B final_adder.U$$135/X final_adder.U$$133/X
+ VGND VGND VPWR VPWR final_adder.U$$261/X sky130_fd_sc_hd__a21o_1
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$100 U$$98/B1 U$$98/A2 U$$924/A1 U$$98/B2 VGND VGND VPWR VPWR U$$101/A sky130_fd_sc_hd__a22o_1
XU$$3939 U$$3939/A U$$3961/B VGND VGND VPWR VPWR U$$3939/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$272 final_adder.U$$274/B final_adder.U$$272/B VGND VGND VPWR VPWR
+ final_adder.U$$398/B sky130_fd_sc_hd__and2_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$111 U$$111/A U$$121/B VGND VGND VPWR VPWR U$$111/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$283 final_adder.U$$282/B final_adder.U$$157/X final_adder.U$$155/X
+ VGND VGND VPWR VPWR final_adder.U$$283/X sky130_fd_sc_hd__a21o_1
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$122 U$$805/B1 U$$98/A2 U$$672/A1 U$$98/B2 VGND VGND VPWR VPWR U$$123/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_32_3 dadda_fa_3_32_3/A dadda_fa_3_32_3/B dadda_fa_3_32_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_33_1/B dadda_fa_4_32_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_73_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$294 final_adder.U$$296/B final_adder.U$$294/B VGND VGND VPWR VPWR
+ final_adder.U$$420/B sky130_fd_sc_hd__and2_1
XU$$133 U$$133/A U$$3/A VGND VGND VPWR VPWR U$$133/X sky130_fd_sc_hd__xor2_1
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$144 U$$144/A U$$180/B VGND VGND VPWR VPWR U$$144/X sky130_fd_sc_hd__xor2_1
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$155 U$$18/A1 U$$179/A2 U$$20/A1 U$$179/B2 VGND VGND VPWR VPWR U$$156/A sky130_fd_sc_hd__a22o_1
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_25_2 U$$1520/X U$$1653/X input174/X VGND VGND VPWR VPWR dadda_fa_4_26_1/A
+ dadda_fa_4_25_2/B sky130_fd_sc_hd__fa_1
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$166 U$$166/A U$$182/B VGND VGND VPWR VPWR U$$166/X sky130_fd_sc_hd__xor2_1
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$177 U$$314/A1 U$$213/A2 U$$42/A1 U$$213/B2 VGND VGND VPWR VPWR U$$178/A sky130_fd_sc_hd__a22o_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$188 U$$188/A U$$220/B VGND VGND VPWR VPWR U$$188/X sky130_fd_sc_hd__xor2_1
XU$$199 U$$62/A1 U$$229/A2 U$$64/A1 U$$229/B2 VGND VGND VPWR VPWR U$$200/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_18_1 U$$442/X U$$575/X U$$708/X VGND VGND VPWR VPWR dadda_fa_4_19_1/B
+ dadda_fa_4_18_2/B sky130_fd_sc_hd__fa_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_396_ _397_/CLK _396_/D VGND VGND VPWR VPWR _396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_77_5 dadda_fa_2_77_5/A dadda_fa_2_77_5/B dadda_fa_2_77_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_2/A dadda_fa_4_77_0/A sky130_fd_sc_hd__fa_2
XFILLER_95_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_886 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_107_1 dadda_fa_5_107_1/A dadda_fa_5_107_1/B dadda_fa_5_107_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_108_0/B dadda_fa_7_107_0/A sky130_fd_sc_hd__fa_1
XFILLER_160_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_858 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout402 U$$807/A2 VGND VGND VPWR VPWR U$$809/A2 sky130_fd_sc_hd__buf_4
XFILLER_59_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout413 U$$642/A2 VGND VGND VPWR VPWR U$$638/A2 sky130_fd_sc_hd__buf_4
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout424 U$$4251/X VGND VGND VPWR VPWR U$$4309/A2 sky130_fd_sc_hd__buf_2
Xdadda_fa_1_72_4 U$$3609/X U$$3742/X U$$3875/X VGND VGND VPWR VPWR dadda_fa_2_73_1/CIN
+ dadda_fa_2_72_4/CIN sky130_fd_sc_hd__fa_1
Xfanout435 U$$4114/X VGND VGND VPWR VPWR U$$4244/A2 sky130_fd_sc_hd__buf_6
Xfanout446 U$$74/A2 VGND VGND VPWR VPWR U$$80/A2 sky130_fd_sc_hd__buf_2
XFILLER_141_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout457 U$$4057/A2 VGND VGND VPWR VPWR U$$4093/A2 sky130_fd_sc_hd__buf_2
Xfanout468 U$$3777/A2 VGND VGND VPWR VPWR U$$3757/A2 sky130_fd_sc_hd__buf_4
XFILLER_171_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_65_3 U$$3728/X U$$3861/X U$$3994/X VGND VGND VPWR VPWR dadda_fa_2_66_1/B
+ dadda_fa_2_65_4/B sky130_fd_sc_hd__fa_1
XFILLER_150_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout479 U$$3658/A2 VGND VGND VPWR VPWR U$$3656/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_86_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_42_2 dadda_fa_4_42_2/A dadda_fa_4_42_2/B dadda_fa_4_42_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_43_0/CIN dadda_fa_5_42_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_58_2 U$$2384/X U$$2517/X U$$2650/X VGND VGND VPWR VPWR dadda_fa_2_59_1/A
+ dadda_fa_2_58_4/A sky130_fd_sc_hd__fa_1
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_35_1 dadda_fa_4_35_1/A dadda_fa_4_35_1/B dadda_fa_4_35_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_36_0/B dadda_fa_5_35_1/B sky130_fd_sc_hd__fa_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_12_0 dadda_fa_7_12_0/A dadda_fa_7_12_0/B dadda_fa_7_12_0/CIN VGND VGND
+ VPWR VPWR _309_/D _180_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_28_0 dadda_fa_4_28_0/A dadda_fa_4_28_0/B dadda_fa_4_28_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_29_0/A dadda_fa_5_28_1/A sky130_fd_sc_hd__fa_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_250_ _391_/CLK _250_/D VGND VGND VPWR VPWR _250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_181_ _344_/CLK _181_/D VGND VGND VPWR VPWR _181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_61_4 U$$1725/X U$$1858/X VGND VGND VPWR VPWR dadda_fa_1_62_7/A dadda_fa_2_61_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_123_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4404 U$$4404/A1 U$$4388/X U$$981/A1 U$$4508/B2 VGND VGND VPWR VPWR U$$4405/A sky130_fd_sc_hd__a22o_1
XU$$4415 U$$4415/A U$$4415/B VGND VGND VPWR VPWR U$$4415/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_60_2 U$$925/X U$$1058/X U$$1191/X VGND VGND VPWR VPWR dadda_fa_1_61_6/CIN
+ dadda_fa_1_60_8/B sky130_fd_sc_hd__fa_1
XU$$4426 U$$4426/A1 U$$4388/X U$$4428/A1 U$$4428/B2 VGND VGND VPWR VPWR U$$4427/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout980 U$$215/B1 VGND VGND VPWR VPWR U$$80/A1 sky130_fd_sc_hd__buf_4
XU$$4437 U$$4437/A U$$4437/B VGND VGND VPWR VPWR U$$4437/X sky130_fd_sc_hd__xor2_1
Xfanout991 U$$4462/A1 VGND VGND VPWR VPWR U$$4460/B1 sky130_fd_sc_hd__buf_4
XFILLER_37_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3703 U$$3701/Y input50/X U$$3699/A U$$3702/X U$$3699/Y VGND VGND VPWR VPWR U$$3703/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_92_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4448 input85/X U$$4388/X U$$4450/A1 U$$4458/B2 VGND VGND VPWR VPWR U$$4449/A sky130_fd_sc_hd__a22o_1
XU$$3714 U$$3714/A U$$3734/B VGND VGND VPWR VPWR U$$3714/X sky130_fd_sc_hd__xor2_1
XU$$4459 U$$4459/A U$$4459/B VGND VGND VPWR VPWR U$$4459/X sky130_fd_sc_hd__xor2_1
XFILLER_161_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3725 U$$3999/A1 U$$3757/A2 U$$3999/B1 U$$3757/B2 VGND VGND VPWR VPWR U$$3726/A
+ sky130_fd_sc_hd__a22o_1
XU$$3736 U$$3736/A U$$3740/B VGND VGND VPWR VPWR U$$3736/X sky130_fd_sc_hd__xor2_1
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3747 U$$3884/A1 U$$3791/A2 U$$4434/A1 U$$3791/B2 VGND VGND VPWR VPWR U$$3748/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3758 U$$3758/A U$$3774/B VGND VGND VPWR VPWR U$$3758/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_30_0 U$$1929/X U$$2062/X U$$2096/B VGND VGND VPWR VPWR dadda_fa_4_31_0/B
+ dadda_fa_4_30_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3769 U$$4043/A1 U$$3773/A2 U$$4043/B1 U$$3773/B2 VGND VGND VPWR VPWR U$$3770/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_379_ _397_/CLK _379_/D VGND VGND VPWR VPWR _379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_82_3 dadda_fa_2_82_3/A dadda_fa_2_82_3/B dadda_fa_2_82_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_1/B dadda_fa_3_82_3/B sky130_fd_sc_hd__fa_1
XFILLER_130_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_75_2 dadda_fa_2_75_2/A dadda_fa_2_75_2/B dadda_fa_2_75_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_1/A dadda_fa_3_75_3/A sky130_fd_sc_hd__fa_1
XFILLER_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_52_1 dadda_fa_5_52_1/A dadda_fa_5_52_1/B dadda_fa_5_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_53_0/B dadda_fa_7_52_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_68_1 dadda_fa_2_68_1/A dadda_fa_2_68_1/B dadda_fa_2_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_0/CIN dadda_fa_3_68_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_45_0 dadda_fa_5_45_0/A dadda_fa_5_45_0/B dadda_fa_5_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_46_0/A dadda_fa_6_45_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1011 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1208 U$$4416/B1 VGND VGND VPWR VPWR U$$3048/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_133_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1219 U$$987/B1 VGND VGND VPWR VPWR U$$2631/B1 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_1_70_1 U$$2674/X U$$2807/X U$$2940/X VGND VGND VPWR VPWR dadda_fa_2_71_0/CIN
+ dadda_fa_2_70_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_8_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_63_0 U$$2394/X U$$2527/X U$$2660/X VGND VGND VPWR VPWR dadda_fa_2_64_0/B
+ dadda_fa_2_63_3/B sky130_fd_sc_hd__fa_1
XFILLER_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2309 U$$2309/A U$$2329/A VGND VGND VPWR VPWR U$$2309/X sky130_fd_sc_hd__xor2_1
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1608 U$$1608/A U$$1608/B VGND VGND VPWR VPWR U$$1608/X sky130_fd_sc_hd__xor2_1
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1619 U$$4220/B1 U$$1625/A2 U$$4361/A1 U$$1625/B2 VGND VGND VPWR VPWR U$$1620/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_302_ _319_/CLK _302_/D VGND VGND VPWR VPWR _302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_233_ _364_/CLK _233_/D VGND VGND VPWR VPWR _233_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_92_2 dadda_fa_3_92_2/A dadda_fa_3_92_2/B dadda_fa_3_92_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_1/A dadda_fa_4_92_2/B sky130_fd_sc_hd__fa_1
XFILLER_171_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_85_1 dadda_fa_3_85_1/A dadda_fa_3_85_1/B dadda_fa_3_85_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_0/CIN dadda_fa_4_85_2/A sky130_fd_sc_hd__fa_1
XFILLER_124_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_62_0 dadda_fa_6_62_0/A dadda_fa_6_62_0/B dadda_fa_6_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_63_0/B dadda_fa_7_62_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_78_0 dadda_fa_3_78_0/A dadda_fa_3_78_0/B dadda_fa_3_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_0/B dadda_fa_4_78_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_112_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_0_52_0 U$$111/X U$$244/X VGND VGND VPWR VPWR dadda_fa_1_53_8/CIN dadda_fa_2_52_0/A
+ sky130_fd_sc_hd__ha_1
Xfanout1720 U$$922/B1 VGND VGND VPWR VPWR U$$2840/B1 sky130_fd_sc_hd__buf_4
Xfanout1731 input105/X VGND VGND VPWR VPWR U$$783/B1 sky130_fd_sc_hd__clkbuf_2
Xfanout1742 U$$3249/A1 VGND VGND VPWR VPWR U$$4482/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1753 U$$3243/B1 VGND VGND VPWR VPWR U$$94/A1 sky130_fd_sc_hd__buf_4
XU$$4201 U$$4201/A U$$4227/B VGND VGND VPWR VPWR U$$4201/X sky130_fd_sc_hd__xor2_1
Xfanout1764 U$$3243/A1 VGND VGND VPWR VPWR U$$3106/A1 sky130_fd_sc_hd__buf_4
XU$$4212 U$$4349/A1 U$$4224/A2 U$$4349/B1 U$$4224/B2 VGND VGND VPWR VPWR U$$4213/A
+ sky130_fd_sc_hd__a22o_1
XU$$4223 U$$4223/A U$$4227/B VGND VGND VPWR VPWR U$$4223/X sky130_fd_sc_hd__xor2_1
Xfanout1775 U$$912/A1 VGND VGND VPWR VPWR U$$773/B1 sky130_fd_sc_hd__buf_6
XU$$4234 U$$4234/A1 U$$4240/A2 U$$4234/B1 U$$4240/B2 VGND VGND VPWR VPWR U$$4235/A
+ sky130_fd_sc_hd__a22o_1
XU$$3500 U$$3500/A U$$3506/B VGND VGND VPWR VPWR U$$3500/X sky130_fd_sc_hd__xor2_1
XU$$4245 U$$4245/A U$$4247/A VGND VGND VPWR VPWR U$$4245/X sky130_fd_sc_hd__xor2_1
XU$$4256 U$$4256/A U$$4292/B VGND VGND VPWR VPWR U$$4256/X sky130_fd_sc_hd__xor2_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3511 U$$4470/A1 U$$3511/A2 U$$3650/A1 U$$3511/B2 VGND VGND VPWR VPWR U$$3512/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4267 U$$4404/A1 U$$4289/A2 U$$981/A1 U$$4289/B2 VGND VGND VPWR VPWR U$$4268/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_114_1 U$$4491/X input145/X dadda_fa_4_114_1/CIN VGND VGND VPWR VPWR dadda_fa_5_115_0/B
+ dadda_fa_5_114_1/B sky130_fd_sc_hd__fa_1
XU$$3522 U$$3522/A U$$3524/B VGND VGND VPWR VPWR U$$3522/X sky130_fd_sc_hd__xor2_1
XFILLER_37_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3533 U$$4081/A1 U$$3559/A2 U$$4081/B1 U$$3559/B2 VGND VGND VPWR VPWR U$$3534/A
+ sky130_fd_sc_hd__a22o_1
XU$$4278 U$$4278/A U$$4322/B VGND VGND VPWR VPWR U$$4278/X sky130_fd_sc_hd__xor2_1
XU$$4289 U$$4424/B1 U$$4289/A2 U$$4291/A1 U$$4289/B2 VGND VGND VPWR VPWR U$$4290/A
+ sky130_fd_sc_hd__a22o_1
XU$$3544 U$$3544/A U$$3561/A VGND VGND VPWR VPWR U$$3544/X sky130_fd_sc_hd__xor2_1
XFILLER_34_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2810 U$$479/B1 U$$2856/A2 U$$346/A1 U$$2856/B2 VGND VGND VPWR VPWR U$$2811/A sky130_fd_sc_hd__a22o_1
XU$$3555 U$$4375/B1 U$$3557/A2 U$$4240/B1 U$$3557/B2 VGND VGND VPWR VPWR U$$3556/A
+ sky130_fd_sc_hd__a22o_1
XU$$3566 U$$3564/Y input48/X U$$3562/A U$$3565/X U$$3562/Y VGND VGND VPWR VPWR U$$3566/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_74_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_107_0 dadda_fa_4_107_0/A dadda_fa_4_107_0/B dadda_fa_4_107_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_108_0/A dadda_fa_5_107_1/A sky130_fd_sc_hd__fa_1
XU$$2821 U$$2821/A U$$2871/B VGND VGND VPWR VPWR U$$2821/X sky130_fd_sc_hd__xor2_1
XU$$2832 U$$3106/A1 U$$2840/A2 U$$3106/B1 U$$2840/B2 VGND VGND VPWR VPWR U$$2833/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3577 U$$3577/A U$$3615/B VGND VGND VPWR VPWR U$$3577/X sky130_fd_sc_hd__xor2_1
XU$$2843 U$$2843/A U$$2877/A VGND VGND VPWR VPWR U$$2843/X sky130_fd_sc_hd__xor2_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3588 U$$3999/A1 U$$3604/A2 U$$3999/B1 U$$3604/B2 VGND VGND VPWR VPWR U$$3589/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3599 U$$3599/A U$$3601/B VGND VGND VPWR VPWR U$$3599/X sky130_fd_sc_hd__xor2_1
XU$$2854 U$$3948/B1 U$$2872/A2 U$$3815/A1 U$$2872/B2 VGND VGND VPWR VPWR U$$2855/A
+ sky130_fd_sc_hd__a22o_1
XU$$2865 U$$2865/A U$$2871/B VGND VGND VPWR VPWR U$$2865/X sky130_fd_sc_hd__xor2_1
XFILLER_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2876 U$$2876/A VGND VGND VPWR VPWR U$$2876/Y sky130_fd_sc_hd__inv_1
XU$$2887 U$$3022/B1 U$$2929/A2 U$$2887/B1 U$$2929/B2 VGND VGND VPWR VPWR U$$2888/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2898 U$$2898/A U$$2938/B VGND VGND VPWR VPWR U$$2898/X sky130_fd_sc_hd__xor2_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_80_0 input235/X dadda_fa_2_80_0/B dadda_fa_2_80_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_81_0/B dadda_fa_3_80_2/B sky130_fd_sc_hd__fa_1
XFILLER_143_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_50_8 U$$3299/X U$$3432/X VGND VGND VPWR VPWR dadda_fa_2_51_3/A dadda_fa_3_50_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$805 final_adder.U$$772/A final_adder.U$$725/X final_adder.U$$693/X
+ VGND VGND VPWR VPWR final_adder.U$$805/X sky130_fd_sc_hd__a21o_1
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$827 final_adder.U$$794/A final_adder.U$$503/X final_adder.U$$715/X
+ VGND VGND VPWR VPWR final_adder.U$$827/X sky130_fd_sc_hd__a21o_1
XFILLER_69_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$849 final_adder.U$$752/X final_adder.U$$817/X final_adder.U$$753/X
+ VGND VGND VPWR VPWR final_adder.U$$849/X sky130_fd_sc_hd__a21o_2
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_95_0 dadda_fa_4_95_0/A dadda_fa_4_95_0/B dadda_fa_4_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_96_0/A dadda_fa_5_95_1/A sky130_fd_sc_hd__fa_1
XFILLER_152_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_109_2 U$$3949/X U$$4082/X U$$4215/X VGND VGND VPWR VPWR dadda_fa_4_110_1/A
+ dadda_fa_4_109_2/B sky130_fd_sc_hd__fa_1
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput380 output380/A VGND VGND VPWR VPWR o[96] sky130_fd_sc_hd__buf_2
XFILLER_105_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1005 fanout1011/X VGND VGND VPWR VPWR U$$74/A1 sky130_fd_sc_hd__buf_4
XFILLER_160_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1016 U$$4182/A1 VGND VGND VPWR VPWR U$$3495/B1 sky130_fd_sc_hd__buf_6
Xfanout1027 U$$1221/B VGND VGND VPWR VPWR U$$1227/B sky130_fd_sc_hd__buf_6
XFILLER_86_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1038 U$$4452/A1 VGND VGND VPWR VPWR U$$68/A1 sky130_fd_sc_hd__buf_4
XFILLER_120_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1049 U$$697/A1 VGND VGND VPWR VPWR U$$12/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2106 U$$2106/A U$$2106/B VGND VGND VPWR VPWR U$$2106/X sky130_fd_sc_hd__xor2_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2117 U$$745/B1 U$$2147/A2 U$$612/A1 U$$2147/B2 VGND VGND VPWR VPWR U$$2118/A sky130_fd_sc_hd__a22o_1
XU$$2128 U$$2128/A U$$2130/B VGND VGND VPWR VPWR U$$2128/X sky130_fd_sc_hd__xor2_1
XFILLER_28_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2139 U$$632/A1 U$$2139/A2 U$$86/A1 U$$2139/B2 VGND VGND VPWR VPWR U$$2140/A sky130_fd_sc_hd__a22o_1
XFILLER_74_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1405 U$$1405/A U$$1415/B VGND VGND VPWR VPWR U$$1405/X sky130_fd_sc_hd__xor2_1
XU$$1416 U$$868/A1 U$$1432/A2 U$$596/A1 U$$1432/B2 VGND VGND VPWR VPWR U$$1417/A sky130_fd_sc_hd__a22o_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1427 U$$1427/A U$$1427/B VGND VGND VPWR VPWR U$$1427/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1438 U$$616/A1 U$$1452/A2 U$$481/A1 U$$1452/B2 VGND VGND VPWR VPWR U$$1439/A sky130_fd_sc_hd__a22o_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1449 U$$1449/A U$$1449/B VGND VGND VPWR VPWR U$$1449/X sky130_fd_sc_hd__xor2_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_216_ _345_/CLK _216_/D VGND VGND VPWR VPWR _216_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1550 input123/X VGND VGND VPWR VPWR U$$4516/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1561 U$$3692/A1 VGND VGND VPWR VPWR U$$3418/A1 sky130_fd_sc_hd__buf_4
XFILLER_38_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1572 input121/X VGND VGND VPWR VPWR U$$3825/B1 sky130_fd_sc_hd__clkbuf_2
XU$$4020 U$$4020/A U$$4110/A VGND VGND VPWR VPWR U$$4020/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_52_4 dadda_fa_2_52_4/A dadda_fa_2_52_4/B dadda_fa_2_52_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_1/CIN dadda_fa_3_52_3/CIN sky130_fd_sc_hd__fa_1
XU$$4031 U$$4440/B1 U$$4045/A2 U$$4307/A1 U$$4045/B2 VGND VGND VPWR VPWR U$$4032/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1583 U$$127/B VGND VGND VPWR VPWR U$$87/B sky130_fd_sc_hd__buf_6
XFILLER_120_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4042 U$$4042/A U$$4110/A VGND VGND VPWR VPWR U$$4042/X sky130_fd_sc_hd__xor2_1
Xfanout1594 input119/X VGND VGND VPWR VPWR U$$811/A1 sky130_fd_sc_hd__clkbuf_8
XU$$4053 U$$215/B1 U$$4057/A2 U$$80/B1 U$$4057/B2 VGND VGND VPWR VPWR U$$4054/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_45_3 dadda_fa_2_45_3/A dadda_fa_2_45_3/B dadda_fa_2_45_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_46_1/B dadda_fa_3_45_3/B sky130_fd_sc_hd__fa_1
XU$$4064 U$$4064/A U$$4082/B VGND VGND VPWR VPWR U$$4064/X sky130_fd_sc_hd__xor2_1
XU$$3330 U$$4426/A1 U$$3338/A2 U$$4428/A1 U$$3338/B2 VGND VGND VPWR VPWR U$$3331/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4075 U$$4484/B1 U$$4081/A2 U$$4488/A1 U$$4081/B2 VGND VGND VPWR VPWR U$$4076/A
+ sky130_fd_sc_hd__a22o_1
XU$$3341 U$$3341/A U$$3341/B VGND VGND VPWR VPWR U$$3341/X sky130_fd_sc_hd__xor2_1
XU$$4086 U$$4086/A U$$4098/B VGND VGND VPWR VPWR U$$4086/X sky130_fd_sc_hd__xor2_1
XU$$3352 U$$4446/B1 U$$3422/A2 U$$4450/A1 U$$3422/B2 VGND VGND VPWR VPWR U$$3353/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_38_2 U$$1945/X U$$2078/X U$$2211/X VGND VGND VPWR VPWR dadda_fa_3_39_1/A
+ dadda_fa_3_38_3/A sky130_fd_sc_hd__fa_1
XU$$4097 U$$4234/A1 U$$4107/A2 U$$4508/B1 U$$4107/B2 VGND VGND VPWR VPWR U$$4098/A
+ sky130_fd_sc_hd__a22o_1
XU$$3363 U$$3363/A U$$3373/B VGND VGND VPWR VPWR U$$3363/X sky130_fd_sc_hd__xor2_1
XU$$3374 U$$3509/B1 U$$3378/A2 U$$3376/A1 U$$3378/B2 VGND VGND VPWR VPWR U$$3375/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_15_1 dadda_fa_5_15_1/A dadda_fa_5_15_1/B dadda_fa_5_15_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_16_0/B dadda_fa_7_15_0/A sky130_fd_sc_hd__fa_2
XU$$3385 U$$3385/A U$$3424/A VGND VGND VPWR VPWR U$$3385/X sky130_fd_sc_hd__xor2_1
XU$$2640 U$$2640/A U$$2678/B VGND VGND VPWR VPWR U$$2640/X sky130_fd_sc_hd__xor2_1
XU$$3396 U$$4081/A1 U$$3416/A2 U$$4081/B1 U$$3416/B2 VGND VGND VPWR VPWR U$$3397/A
+ sky130_fd_sc_hd__a22o_1
XU$$2651 U$$2925/A1 U$$2667/A2 U$$3338/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2652/A
+ sky130_fd_sc_hd__a22o_1
XU$$2662 U$$2662/A U$$2662/B VGND VGND VPWR VPWR U$$2662/X sky130_fd_sc_hd__xor2_1
XFILLER_62_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2673 U$$4454/A1 U$$2707/A2 U$$3495/B1 U$$2707/B2 VGND VGND VPWR VPWR U$$2674/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2684 U$$2684/A U$$2739/A VGND VGND VPWR VPWR U$$2684/X sky130_fd_sc_hd__xor2_1
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2695 U$$3106/A1 U$$2707/A2 U$$3106/B1 U$$2707/B2 VGND VGND VPWR VPWR U$$2696/A
+ sky130_fd_sc_hd__a22o_1
XU$$1950 U$$991/A1 U$$2006/A2 U$$854/B1 U$$2006/B2 VGND VGND VPWR VPWR U$$1951/A sky130_fd_sc_hd__a22o_1
XFILLER_22_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1961 U$$1961/A U$$1963/B VGND VGND VPWR VPWR U$$1961/X sky130_fd_sc_hd__xor2_1
XU$$1972 U$$739/A1 U$$1980/A2 U$$741/A1 U$$1980/B2 VGND VGND VPWR VPWR U$$1973/A sky130_fd_sc_hd__a22o_1
XU$$1983 U$$1983/A U$$2015/B VGND VGND VPWR VPWR U$$1983/X sky130_fd_sc_hd__xor2_1
XU$$1994 U$$3636/B1 U$$2046/A2 U$$3638/B1 U$$2046/B2 VGND VGND VPWR VPWR U$$1995/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput108 b[49] VGND VGND VPWR VPWR input108/X sky130_fd_sc_hd__clkbuf_1
Xinput119 b[59] VGND VGND VPWR VPWR input119/X sky130_fd_sc_hd__buf_2
XFILLER_69_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$602 final_adder.U$$610/B final_adder.U$$602/B VGND VGND VPWR VPWR
+ final_adder.U$$706/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$613 final_adder.U$$612/B final_adder.U$$497/X final_adder.U$$489/X
+ VGND VGND VPWR VPWR final_adder.U$$613/X sky130_fd_sc_hd__a21o_1
XFILLER_111_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$635 final_adder.U$$634/B final_adder.U$$531/X final_adder.U$$515/X
+ VGND VGND VPWR VPWR final_adder.U$$635/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$646 final_adder.U$$662/B final_adder.U$$646/B VGND VGND VPWR VPWR
+ final_adder.U$$758/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$657 final_adder.U$$656/B final_adder.U$$553/X final_adder.U$$537/X
+ VGND VGND VPWR VPWR final_adder.U$$657/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$668 final_adder.U$$684/B final_adder.U$$668/B VGND VGND VPWR VPWR
+ final_adder.U$$780/B sky130_fd_sc_hd__and2_1
XU$$507 U$$918/A1 U$$545/A2 U$$920/A1 U$$545/B2 VGND VGND VPWR VPWR U$$508/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$679 final_adder.U$$678/B final_adder.U$$575/X final_adder.U$$559/X
+ VGND VGND VPWR VPWR final_adder.U$$679/X sky130_fd_sc_hd__a21o_1
XFILLER_38_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$518 U$$518/A U$$522/B VGND VGND VPWR VPWR U$$518/X sky130_fd_sc_hd__xor2_1
XU$$529 U$$803/A1 U$$539/A2 U$$805/A1 U$$539/B2 VGND VGND VPWR VPWR U$$530/A sky130_fd_sc_hd__a22o_1
XFILLER_38_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_40_2 U$$885/X U$$1018/X U$$1151/X VGND VGND VPWR VPWR dadda_fa_2_41_4/B
+ dadda_fa_2_40_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$90 U$$90/A1 U$$96/A2 U$$92/A1 U$$96/B2 VGND VGND VPWR VPWR U$$91/A sky130_fd_sc_hd__a22o_1
XFILLER_25_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_10_0 U$$27/X U$$160/X U$$293/X VGND VGND VPWR VPWR dadda_fa_5_11_0/CIN
+ dadda_fa_5_10_1/B sky130_fd_sc_hd__fa_1
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_114_0 dadda_fa_3_114_0/A U$$3560/X U$$3693/X VGND VGND VPWR VPWR dadda_fa_4_115_2/A
+ dadda_fa_4_114_2/B sky130_fd_sc_hd__fa_1
XFILLER_122_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_62_3 dadda_fa_3_62_3/A dadda_fa_3_62_3/B dadda_fa_3_62_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_1/B dadda_fa_4_62_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_55_2 dadda_fa_3_55_2/A dadda_fa_3_55_2/B dadda_fa_3_55_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_1/A dadda_fa_4_55_2/B sky130_fd_sc_hd__fa_1
XFILLER_48_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_48_1 dadda_fa_3_48_1/A dadda_fa_3_48_1/B dadda_fa_3_48_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_0/CIN dadda_fa_4_48_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_25_0 dadda_fa_6_25_0/A dadda_fa_6_25_0/B dadda_fa_6_25_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_26_0/B dadda_fa_7_25_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_62_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1202 U$$928/A1 U$$1202/A2 U$$930/A1 U$$1202/B2 VGND VGND VPWR VPWR U$$1203/A sky130_fd_sc_hd__a22o_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1213 U$$1213/A U$$1227/B VGND VGND VPWR VPWR U$$1213/X sky130_fd_sc_hd__xor2_1
XU$$1224 U$$539/A1 U$$1226/A2 U$$678/A1 U$$1226/B2 VGND VGND VPWR VPWR U$$1225/A sky130_fd_sc_hd__a22o_1
XU$$1235 U$$1370/A VGND VGND VPWR VPWR U$$1235/Y sky130_fd_sc_hd__inv_1
XFILLER_90_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1246 U$$1246/A U$$1282/B VGND VGND VPWR VPWR U$$1246/X sky130_fd_sc_hd__xor2_1
XU$$1257 U$$983/A1 U$$1295/A2 U$$983/B1 U$$1295/B2 VGND VGND VPWR VPWR U$$1258/A sky130_fd_sc_hd__a22o_1
XU$$1268 U$$1268/A U$$1282/B VGND VGND VPWR VPWR U$$1268/X sky130_fd_sc_hd__xor2_1
XU$$1279 U$$183/A1 U$$1311/A2 U$$48/A1 U$$1311/B2 VGND VGND VPWR VPWR U$$1280/A sky130_fd_sc_hd__a22o_1
XFILLER_129_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1040 final_adder.U$$238/A final_adder.U$$619/X VGND VGND VPWR VPWR
+ output292/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1051 final_adder.U$$228/B final_adder.U$$999/X VGND VGND VPWR VPWR
+ output304/A sky130_fd_sc_hd__xor2_1
XFILLER_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1062 final_adder.U$$216/A final_adder.U$$829/X VGND VGND VPWR VPWR
+ output316/A sky130_fd_sc_hd__xor2_1
XFILLER_171_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1073 final_adder.U$$206/B final_adder.U$$977/X VGND VGND VPWR VPWR
+ output328/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1084 final_adder.U$$194/A final_adder.U$$807/X VGND VGND VPWR VPWR
+ output341/A sky130_fd_sc_hd__xor2_1
XFILLER_116_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1095 final_adder.U$$184/B final_adder.U$$955/X VGND VGND VPWR VPWR
+ output353/A sky130_fd_sc_hd__xor2_1
XFILLER_98_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout809 U$$2733/B2 VGND VGND VPWR VPWR U$$2737/B2 sky130_fd_sc_hd__buf_4
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_50_1 dadda_fa_2_50_1/A dadda_fa_2_50_1/B dadda_fa_2_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_0/CIN dadda_fa_3_50_2/CIN sky130_fd_sc_hd__fa_1
Xfanout1380 U$$2986/B VGND VGND VPWR VPWR U$$3013/A sky130_fd_sc_hd__buf_2
Xfanout1391 input36/X VGND VGND VPWR VPWR fanout1391/X sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_2_43_0 U$$1955/X U$$2088/X U$$2221/X VGND VGND VPWR VPWR dadda_fa_3_44_0/B
+ dadda_fa_3_43_2/B sky130_fd_sc_hd__fa_1
XFILLER_81_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$545_1908 VGND VGND VPWR VPWR U$$545_1908/HI U$$545/B1 sky130_fd_sc_hd__conb_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3160 U$$3160/A U$$3196/B VGND VGND VPWR VPWR U$$3160/X sky130_fd_sc_hd__xor2_1
XU$$3171 U$$979/A1 U$$3257/A2 U$$979/B1 U$$3257/B2 VGND VGND VPWR VPWR U$$3172/A sky130_fd_sc_hd__a22o_1
XFILLER_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3182 U$$3182/A U$$3210/B VGND VGND VPWR VPWR U$$3182/X sky130_fd_sc_hd__xor2_1
XU$$3193 U$$4426/A1 U$$3199/A2 U$$4428/A1 U$$3199/B2 VGND VGND VPWR VPWR U$$3194/A
+ sky130_fd_sc_hd__a22o_1
XU$$2470 U$$2468/Y input30/X U$$2466/A U$$2469/X U$$2466/Y VGND VGND VPWR VPWR U$$2470/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_50_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2481 U$$2481/A U$$2541/B VGND VGND VPWR VPWR U$$2481/X sky130_fd_sc_hd__xor2_1
XU$$2492 U$$2629/A1 U$$2532/A2 U$$2631/A1 U$$2532/B2 VGND VGND VPWR VPWR U$$2493/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1780 U$$1781/A VGND VGND VPWR VPWR U$$1780/Y sky130_fd_sc_hd__inv_1
XU$$1791 U$$3022/B1 U$$1829/A2 U$$2887/B1 U$$1829/B2 VGND VGND VPWR VPWR U$$1792/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput90 b[32] VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_72_2 dadda_fa_4_72_2/A dadda_fa_4_72_2/B dadda_fa_4_72_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_73_0/CIN dadda_fa_5_72_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_162_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_88_2 U$$2444/X U$$2577/X U$$2710/X VGND VGND VPWR VPWR dadda_fa_2_89_4/A
+ dadda_fa_2_88_5/B sky130_fd_sc_hd__fa_1
Xdadda_fa_4_65_1 dadda_fa_4_65_1/A dadda_fa_4_65_1/B dadda_fa_4_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_66_0/B dadda_fa_5_65_1/B sky130_fd_sc_hd__fa_1
XFILLER_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_42_0 dadda_fa_7_42_0/A dadda_fa_7_42_0/B dadda_fa_7_42_0/CIN VGND VGND
+ VPWR VPWR _339_/D _210_/D sky130_fd_sc_hd__fa_2
XFILLER_76_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_58_0 dadda_fa_4_58_0/A dadda_fa_4_58_0/B dadda_fa_4_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_59_0/A dadda_fa_5_58_1/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$410 final_adder.U$$414/B final_adder.U$$410/B VGND VGND VPWR VPWR
+ final_adder.U$$534/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$421 final_adder.U$$420/B final_adder.U$$299/X final_adder.U$$295/X
+ VGND VGND VPWR VPWR final_adder.U$$421/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$432 final_adder.U$$436/B final_adder.U$$432/B VGND VGND VPWR VPWR
+ final_adder.U$$556/B sky130_fd_sc_hd__and2_1
XFILLER_123_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$443 final_adder.U$$442/B final_adder.U$$321/X final_adder.U$$317/X
+ VGND VGND VPWR VPWR final_adder.U$$443/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$454 final_adder.U$$458/B final_adder.U$$454/B VGND VGND VPWR VPWR
+ final_adder.U$$578/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$465 final_adder.U$$464/B final_adder.U$$343/X final_adder.U$$339/X
+ VGND VGND VPWR VPWR final_adder.U$$465/X sky130_fd_sc_hd__a21o_1
XU$$304 U$$576/B1 U$$338/A2 U$$443/A1 U$$338/B2 VGND VGND VPWR VPWR U$$305/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$476 final_adder.U$$480/B final_adder.U$$476/B VGND VGND VPWR VPWR
+ final_adder.U$$600/B sky130_fd_sc_hd__and2_1
XFILLER_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$315 U$$315/A U$$341/B VGND VGND VPWR VPWR U$$315/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$487 final_adder.U$$486/B final_adder.U$$365/X final_adder.U$$361/X
+ VGND VGND VPWR VPWR final_adder.U$$487/X sky130_fd_sc_hd__a21o_1
XU$$326 U$$598/B1 U$$362/A2 U$$465/A1 U$$362/B2 VGND VGND VPWR VPWR U$$327/A sky130_fd_sc_hd__a22o_1
XFILLER_83_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$498 final_adder.U$$498/A final_adder.U$$498/B VGND VGND VPWR VPWR
+ final_adder.U$$614/A sky130_fd_sc_hd__and2_1
XU$$337 U$$337/A U$$353/B VGND VGND VPWR VPWR U$$337/X sky130_fd_sc_hd__xor2_1
XFILLER_44_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$348 U$$74/A1 U$$352/A2 U$$74/B1 U$$352/B2 VGND VGND VPWR VPWR U$$349/A sky130_fd_sc_hd__a22o_1
XU$$359 U$$359/A U$$363/B VGND VGND VPWR VPWR U$$359/X sky130_fd_sc_hd__xor2_1
XU$$4505_1900 VGND VGND VPWR VPWR U$$4505_1900/HI U$$4505/B sky130_fd_sc_hd__conb_1
XFILLER_32_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_60_0 dadda_fa_3_60_0/A dadda_fa_3_60_0/B dadda_fa_3_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_0/B dadda_fa_4_60_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_76_0 dadda_fa_0_76_0/A U$$957/X U$$1090/X VGND VGND VPWR VPWR dadda_fa_1_77_8/B
+ dadda_fa_1_76_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_110_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$860 U$$997/A1 U$$898/A2 U$$997/B1 U$$898/B2 VGND VGND VPWR VPWR U$$861/A sky130_fd_sc_hd__a22o_1
XU$$871 U$$871/A U$$875/B VGND VGND VPWR VPWR U$$871/X sky130_fd_sc_hd__xor2_1
XU$$1010 U$$1010/A U$$980/B VGND VGND VPWR VPWR U$$1010/X sky130_fd_sc_hd__xor2_1
XU$$1021 U$$62/A1 U$$997/A2 U$$64/A1 U$$997/B2 VGND VGND VPWR VPWR U$$1022/A sky130_fd_sc_hd__a22o_1
XFILLER_51_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$882 U$$882/A1 U$$904/A2 U$$882/B1 U$$904/B2 VGND VGND VPWR VPWR U$$883/A sky130_fd_sc_hd__a22o_1
XU$$1032 U$$1032/A U$$1062/B VGND VGND VPWR VPWR U$$1032/X sky130_fd_sc_hd__xor2_1
XU$$893 U$$893/A U$$895/B VGND VGND VPWR VPWR U$$893/X sky130_fd_sc_hd__xor2_1
XU$$1043 U$$82/B1 U$$1087/A2 U$$906/B1 U$$1087/B2 VGND VGND VPWR VPWR U$$1044/A sky130_fd_sc_hd__a22o_1
XU$$1054 U$$1054/A U$$1094/B VGND VGND VPWR VPWR U$$1054/X sky130_fd_sc_hd__xor2_1
XU$$1065 U$$928/A1 U$$1075/A2 U$$930/A1 U$$1075/B2 VGND VGND VPWR VPWR U$$1066/A sky130_fd_sc_hd__a22o_1
XU$$1076 U$$1076/A U$$990/B VGND VGND VPWR VPWR U$$1076/X sky130_fd_sc_hd__xor2_1
XFILLER_31_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1087 U$$950/A1 U$$1087/A2 U$$952/A1 U$$1087/B2 VGND VGND VPWR VPWR U$$1088/A sky130_fd_sc_hd__a22o_1
XU$$1098 U$$1233/A VGND VGND VPWR VPWR U$$1098/Y sky130_fd_sc_hd__inv_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_82_1 dadda_fa_5_82_1/A dadda_fa_5_82_1/B dadda_fa_5_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_83_0/B dadda_fa_7_82_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_98_1 U$$2730/X U$$2863/X U$$2996/X VGND VGND VPWR VPWR dadda_fa_3_99_1/A
+ dadda_fa_3_98_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_75_0 dadda_fa_5_75_0/A dadda_fa_5_75_0/B dadda_fa_5_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_76_0/A dadda_fa_6_75_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout606 U$$1720/A2 VGND VGND VPWR VPWR U$$1702/A2 sky130_fd_sc_hd__buf_4
XFILLER_99_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout617 U$$1625/A2 VGND VGND VPWR VPWR U$$1641/A2 sky130_fd_sc_hd__clkbuf_8
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout628 U$$141/X VGND VGND VPWR VPWR U$$253/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_74_8 dadda_fa_1_74_8/A dadda_fa_1_74_8/B dadda_fa_1_74_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_75_3/A dadda_fa_3_74_0/A sky130_fd_sc_hd__fa_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout639 U$$1361/A2 VGND VGND VPWR VPWR U$$1367/A2 sky130_fd_sc_hd__buf_4
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_67_7 dadda_fa_1_67_7/A dadda_fa_1_67_7/B dadda_fa_1_67_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_68_2/CIN dadda_fa_2_67_5/CIN sky130_fd_sc_hd__fa_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_976 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_784 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_93_0 U$$2054/Y U$$2188/X U$$2321/X VGND VGND VPWR VPWR dadda_fa_2_94_5/A
+ dadda_fa_2_93_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3907 U$$3907/A U$$3907/B VGND VGND VPWR VPWR U$$3907/X sky130_fd_sc_hd__xor2_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$240 final_adder.U$$240/A final_adder.U$$240/B VGND VGND VPWR VPWR
+ final_adder.U$$368/B sky130_fd_sc_hd__and2_1
XFILLER_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$251 final_adder.U$$5/SUM final_adder.U$$4/COUT final_adder.U$$5/COUT
+ VGND VGND VPWR VPWR final_adder.U$$251/X sky130_fd_sc_hd__a21o_1
XFILLER_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3918 U$$4464/B1 U$$3948/A2 U$$4331/A1 U$$3948/B2 VGND VGND VPWR VPWR U$$3919/A
+ sky130_fd_sc_hd__a22o_1
XU$$3929 U$$3929/A U$$3949/B VGND VGND VPWR VPWR U$$3929/X sky130_fd_sc_hd__xor2_1
XU$$101 U$$101/A U$$99/B VGND VGND VPWR VPWR U$$101/X sky130_fd_sc_hd__xor2_1
XFILLER_100_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$262 final_adder.U$$264/B final_adder.U$$262/B VGND VGND VPWR VPWR
+ final_adder.U$$388/B sky130_fd_sc_hd__and2_1
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_105_0 dadda_fa_6_105_0/A dadda_fa_6_105_0/B dadda_fa_6_105_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_106_0/B dadda_fa_7_105_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$273 final_adder.U$$272/B final_adder.U$$147/X final_adder.U$$145/X
+ VGND VGND VPWR VPWR final_adder.U$$273/X sky130_fd_sc_hd__a21o_1
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$112 U$$521/B1 U$$120/A2 U$$386/B1 U$$120/B2 VGND VGND VPWR VPWR U$$113/A sky130_fd_sc_hd__a22o_1
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$284 final_adder.U$$286/B final_adder.U$$284/B VGND VGND VPWR VPWR
+ final_adder.U$$410/B sky130_fd_sc_hd__and2_1
XU$$123 U$$123/A U$$127/B VGND VGND VPWR VPWR U$$123/X sky130_fd_sc_hd__xor2_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$295 final_adder.U$$294/B final_adder.U$$169/X final_adder.U$$167/X
+ VGND VGND VPWR VPWR final_adder.U$$295/X sky130_fd_sc_hd__a21o_1
XU$$134 U$$406/B1 U$$98/A2 U$$134/B1 U$$98/B2 VGND VGND VPWR VPWR U$$135/A sky130_fd_sc_hd__a22o_1
XFILLER_45_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$145 U$$965/B1 U$$179/A2 U$$10/A1 U$$179/B2 VGND VGND VPWR VPWR U$$146/A sky130_fd_sc_hd__a22o_1
XFILLER_27_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_25_3 dadda_fa_3_25_3/A dadda_fa_3_25_3/B dadda_fa_3_25_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_26_1/B dadda_fa_4_25_2/CIN sky130_fd_sc_hd__fa_1
XU$$156 U$$156/A U$$180/B VGND VGND VPWR VPWR U$$156/X sky130_fd_sc_hd__xor2_1
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$167 U$$576/B1 U$$207/A2 U$$443/A1 U$$207/B2 VGND VGND VPWR VPWR U$$168/A sky130_fd_sc_hd__a22o_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$178 U$$178/A U$$182/B VGND VGND VPWR VPWR U$$178/X sky130_fd_sc_hd__xor2_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$189 U$$52/A1 U$$219/A2 U$$54/A1 U$$219/B2 VGND VGND VPWR VPWR U$$190/A sky130_fd_sc_hd__a22o_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_395_ _397_/CLK _395_/D VGND VGND VPWR VPWR _395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_92_0 dadda_fa_6_92_0/A dadda_fa_6_92_0/B dadda_fa_6_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_93_0/B dadda_fa_7_92_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_127_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$690 U$$688/B U$$685/A input2/X U$$685/Y VGND VGND VPWR VPWR U$$690/X sky130_fd_sc_hd__a22o_2
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_80_8 U$$4290/X U$$4423/X VGND VGND VPWR VPWR dadda_fa_2_81_3/B dadda_fa_3_80_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_173_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout403 U$$689/X VGND VGND VPWR VPWR U$$807/A2 sky130_fd_sc_hd__buf_4
Xfanout414 U$$642/A2 VGND VGND VPWR VPWR U$$682/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout425 U$$543/A2 VGND VGND VPWR VPWR U$$497/A2 sky130_fd_sc_hd__buf_4
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout436 U$$4190/A2 VGND VGND VPWR VPWR U$$4240/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_72_5 U$$4008/X U$$4141/X U$$4274/X VGND VGND VPWR VPWR dadda_fa_2_73_2/A
+ dadda_fa_2_72_5/A sky130_fd_sc_hd__fa_1
XFILLER_113_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout447 U$$120/A2 VGND VGND VPWR VPWR U$$74/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout458 U$$3977/X VGND VGND VPWR VPWR U$$4057/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_65_4 U$$4127/X U$$4260/X U$$4393/X VGND VGND VPWR VPWR dadda_fa_2_66_1/CIN
+ dadda_fa_2_65_4/CIN sky130_fd_sc_hd__fa_1
Xfanout469 U$$3777/A2 VGND VGND VPWR VPWR U$$3739/A2 sky130_fd_sc_hd__buf_2
XFILLER_101_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_58_3 U$$2783/X U$$2916/X U$$3049/X VGND VGND VPWR VPWR dadda_fa_2_59_1/B
+ dadda_fa_2_58_4/B sky130_fd_sc_hd__fa_1
XFILLER_27_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_35_2 dadda_fa_4_35_2/A dadda_fa_4_35_2/B dadda_fa_4_35_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_36_0/CIN dadda_fa_5_35_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_28_1 dadda_fa_4_28_1/A dadda_fa_4_28_1/B dadda_fa_4_28_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_29_0/B dadda_fa_5_28_1/B sky130_fd_sc_hd__fa_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1006 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_180_ _344_/CLK _180_/D VGND VGND VPWR VPWR _180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4405 U$$4405/A U$$4405/B VGND VGND VPWR VPWR U$$4405/X sky130_fd_sc_hd__xor2_1
Xfanout970 fanout975/X VGND VGND VPWR VPWR U$$3642/B1 sky130_fd_sc_hd__buf_4
XU$$4416 U$$4416/A1 U$$4388/X U$$4416/B1 U$$4506/B2 VGND VGND VPWR VPWR U$$4417/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_0_60_3 U$$1324/X U$$1457/X U$$1590/X VGND VGND VPWR VPWR dadda_fa_1_61_7/A
+ dadda_fa_1_60_8/CIN sky130_fd_sc_hd__fa_1
Xfanout981 fanout984/X VGND VGND VPWR VPWR U$$215/B1 sky130_fd_sc_hd__buf_4
XU$$4427 U$$4427/A U$$4427/B VGND VGND VPWR VPWR U$$4427/X sky130_fd_sc_hd__xor2_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4438 U$$4438/A1 U$$4388/X U$$4440/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4439/A
+ sky130_fd_sc_hd__a22o_1
Xfanout992 fanout993/X VGND VGND VPWR VPWR U$$4462/A1 sky130_fd_sc_hd__buf_4
XFILLER_38_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3704 U$$3702/B U$$3699/A input50/X U$$3699/Y VGND VGND VPWR VPWR U$$3704/X sky130_fd_sc_hd__a22o_4
Xdadda_ha_3_17_1 U$$440/X U$$573/X VGND VGND VPWR VPWR dadda_fa_4_18_1/CIN dadda_ha_3_17_1/SUM
+ sky130_fd_sc_hd__ha_1
XU$$4449 U$$4449/A U$$4449/B VGND VGND VPWR VPWR U$$4449/X sky130_fd_sc_hd__xor2_1
XFILLER_58_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3715 U$$4400/A1 U$$3739/A2 U$$4402/A1 U$$3739/B2 VGND VGND VPWR VPWR U$$3716/A
+ sky130_fd_sc_hd__a22o_1
XU$$3726 U$$3726/A U$$3734/B VGND VGND VPWR VPWR U$$3726/X sky130_fd_sc_hd__xor2_1
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3737 U$$4420/B1 U$$3739/A2 U$$4287/A1 U$$3739/B2 VGND VGND VPWR VPWR U$$3738/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_30_1 input180/X dadda_fa_3_30_1/B dadda_fa_3_30_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_31_0/CIN dadda_fa_4_30_2/A sky130_fd_sc_hd__fa_1
XU$$3748 U$$3748/A U$$3790/B VGND VGND VPWR VPWR U$$3748/X sky130_fd_sc_hd__xor2_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3759 U$$4442/B1 U$$3773/A2 U$$4309/A1 U$$3773/B2 VGND VGND VPWR VPWR U$$3760/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_23_0 U$$319/X U$$452/X U$$585/X VGND VGND VPWR VPWR dadda_fa_4_24_0/B
+ dadda_fa_4_23_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_72_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_378_ _397_/CLK _378_/D VGND VGND VPWR VPWR _378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_82_4 dadda_fa_2_82_4/A dadda_fa_2_82_4/B dadda_fa_2_82_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_1/CIN dadda_fa_3_82_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_75_3 dadda_fa_2_75_3/A dadda_fa_2_75_3/B dadda_fa_2_75_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_1/B dadda_fa_3_75_3/B sky130_fd_sc_hd__fa_1
XFILLER_123_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_68_2 dadda_fa_2_68_2/A dadda_fa_2_68_2/B dadda_fa_2_68_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_1/A dadda_fa_3_68_3/A sky130_fd_sc_hd__fa_1
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_45_1 dadda_fa_5_45_1/A dadda_fa_5_45_1/B dadda_fa_5_45_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_46_0/B dadda_fa_7_45_0/A sky130_fd_sc_hd__fa_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_38_0 dadda_fa_5_38_0/A dadda_fa_5_38_0/B dadda_fa_5_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_39_0/A dadda_fa_6_38_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_37_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1023 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_112_0 dadda_fa_5_112_0/A dadda_fa_5_112_0/B dadda_fa_5_112_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_113_0/A dadda_fa_6_112_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1209 input69/X VGND VGND VPWR VPWR U$$4416/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_70_2 U$$3073/X U$$3206/X U$$3339/X VGND VGND VPWR VPWR dadda_fa_2_71_1/A
+ dadda_fa_2_70_4/A sky130_fd_sc_hd__fa_1
XFILLER_115_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_63_1 U$$2793/X U$$2926/X U$$3059/X VGND VGND VPWR VPWR dadda_fa_2_64_0/CIN
+ dadda_fa_2_63_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_40_0 dadda_fa_4_40_0/A dadda_fa_4_40_0/B dadda_fa_4_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_41_0/A dadda_fa_5_40_1/A sky130_fd_sc_hd__fa_1
XFILLER_75_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_56_0 U$$1183/X U$$1316/X U$$1449/X VGND VGND VPWR VPWR dadda_fa_2_57_0/B
+ dadda_fa_2_56_3/B sky130_fd_sc_hd__fa_1
XFILLER_28_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4385_1837 VGND VGND VPWR VPWR U$$4385_1837/HI U$$4385/A sky130_fd_sc_hd__conb_1
XFILLER_90_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1609 U$$787/A1 U$$1625/A2 U$$787/B1 U$$1625/B2 VGND VGND VPWR VPWR U$$1610/A sky130_fd_sc_hd__a22o_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_301_ _319_/CLK _301_/D VGND VGND VPWR VPWR _301_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_232_ _361_/CLK _232_/D VGND VGND VPWR VPWR _232_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_129_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_92_3 dadda_fa_3_92_3/A dadda_fa_3_92_3/B dadda_fa_3_92_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_1/B dadda_fa_4_92_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_85_2 dadda_fa_3_85_2/A dadda_fa_3_85_2/B dadda_fa_3_85_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_1/A dadda_fa_4_85_2/B sky130_fd_sc_hd__fa_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_78_1 dadda_fa_3_78_1/A dadda_fa_3_78_1/B dadda_fa_3_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_0/CIN dadda_fa_4_78_2/A sky130_fd_sc_hd__fa_1
XFILLER_152_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_55_0 dadda_fa_6_55_0/A dadda_fa_6_55_0/B dadda_fa_6_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_56_0/B dadda_fa_7_55_0/CIN sky130_fd_sc_hd__fa_1
Xfanout1710 U$$2979/B1 VGND VGND VPWR VPWR U$$926/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout1721 input106/X VGND VGND VPWR VPWR U$$922/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout1732 U$$3249/B1 VGND VGND VPWR VPWR U$$4482/B1 sky130_fd_sc_hd__buf_4
XFILLER_78_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1743 input104/X VGND VGND VPWR VPWR U$$3249/A1 sky130_fd_sc_hd__buf_6
Xfanout1754 U$$3243/B1 VGND VGND VPWR VPWR U$$505/A1 sky130_fd_sc_hd__clkbuf_4
XU$$4202 U$$4474/B1 U$$4224/A2 U$$4341/A1 U$$4224/B2 VGND VGND VPWR VPWR U$$4203/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1765 input101/X VGND VGND VPWR VPWR U$$3243/A1 sky130_fd_sc_hd__buf_6
XU$$4213 U$$4213/A U$$4215/B VGND VGND VPWR VPWR U$$4213/X sky130_fd_sc_hd__xor2_1
XU$$4224 U$$4359/B1 U$$4224/A2 U$$4226/A1 U$$4224/B2 VGND VGND VPWR VPWR U$$4225/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1776 U$$3650/B1 VGND VGND VPWR VPWR U$$4198/B1 sky130_fd_sc_hd__buf_4
XU$$4235 U$$4235/A U$$4241/B VGND VGND VPWR VPWR U$$4235/X sky130_fd_sc_hd__xor2_1
XU$$3501 U$$3636/B1 U$$3505/A2 U$$3638/B1 U$$3505/B2 VGND VGND VPWR VPWR U$$3502/A
+ sky130_fd_sc_hd__a22o_1
XU$$4246 U$$4247/A VGND VGND VPWR VPWR U$$4246/Y sky130_fd_sc_hd__inv_1
XU$$4257 U$$4257/A1 U$$4295/A2 U$$4257/B1 U$$4295/B2 VGND VGND VPWR VPWR U$$4258/A
+ sky130_fd_sc_hd__a22o_1
XU$$3512 U$$3512/A U$$3562/A VGND VGND VPWR VPWR U$$3512/X sky130_fd_sc_hd__xor2_1
XU$$4268 U$$4268/A U$$4294/B VGND VGND VPWR VPWR U$$4268/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_114_2 dadda_fa_4_114_2/A dadda_fa_4_114_2/B dadda_ha_3_114_1/SUM VGND
+ VGND VPWR VPWR dadda_fa_5_115_0/CIN dadda_fa_5_114_1/CIN sky130_fd_sc_hd__fa_1
XU$$3523 U$$920/A1 U$$3523/A2 U$$920/B1 U$$3523/B2 VGND VGND VPWR VPWR U$$3524/A sky130_fd_sc_hd__a22o_1
XU$$3534 U$$3534/A U$$3548/B VGND VGND VPWR VPWR U$$3534/X sky130_fd_sc_hd__xor2_1
XU$$4279 U$$4416/A1 U$$4325/A2 U$$4416/B1 U$$4325/B2 VGND VGND VPWR VPWR U$$4280/A
+ sky130_fd_sc_hd__a22o_1
XU$$2800 U$$4442/B1 U$$2804/A2 U$$4309/A1 U$$2804/B2 VGND VGND VPWR VPWR U$$2801/A
+ sky130_fd_sc_hd__a22o_1
XU$$3545 U$$3817/B1 U$$3549/A2 U$$3684/A1 U$$3549/B2 VGND VGND VPWR VPWR U$$3546/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2811 U$$2811/A U$$2811/B VGND VGND VPWR VPWR U$$2811/X sky130_fd_sc_hd__xor2_1
XFILLER_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3556 U$$3556/A U$$3558/B VGND VGND VPWR VPWR U$$3556/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_107_1 dadda_fa_4_107_1/A dadda_fa_4_107_1/B dadda_fa_4_107_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_108_0/B dadda_fa_5_107_1/B sky130_fd_sc_hd__fa_1
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3567 U$$3565/B U$$3562/A input48/X U$$3562/Y VGND VGND VPWR VPWR U$$3567/X sky130_fd_sc_hd__a22o_2
XU$$2822 U$$4466/A1 U$$2874/A2 U$$4468/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2823/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2833 U$$2833/A U$$2841/B VGND VGND VPWR VPWR U$$2833/X sky130_fd_sc_hd__xor2_1
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3578 U$$3713/B1 U$$3656/A2 U$$3580/A1 U$$3656/B2 VGND VGND VPWR VPWR U$$3579/A
+ sky130_fd_sc_hd__a22o_1
XU$$3589 U$$3589/A U$$3601/B VGND VGND VPWR VPWR U$$3589/X sky130_fd_sc_hd__xor2_1
XU$$2844 U$$2979/B1 U$$2844/A2 U$$2844/B1 U$$2844/B2 VGND VGND VPWR VPWR U$$2845/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2855 U$$2855/A U$$2871/B VGND VGND VPWR VPWR U$$2855/X sky130_fd_sc_hd__xor2_1
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2866 U$$3551/A1 U$$2874/A2 U$$3416/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2867/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2877 U$$2877/A VGND VGND VPWR VPWR U$$2877/Y sky130_fd_sc_hd__inv_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2888 U$$2888/A U$$2926/B VGND VGND VPWR VPWR U$$2888/X sky130_fd_sc_hd__xor2_1
XU$$2899 U$$707/A1 U$$2991/A2 U$$709/A1 U$$2991/B2 VGND VGND VPWR VPWR U$$2900/A sky130_fd_sc_hd__a22o_1
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_80_1 dadda_fa_2_80_1/A dadda_fa_2_80_1/B dadda_fa_2_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_0/CIN dadda_fa_3_80_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_73_0 dadda_fa_2_73_0/A dadda_fa_2_73_0/B dadda_fa_2_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_0/B dadda_fa_3_73_2/B sky130_fd_sc_hd__fa_1
XFILLER_170_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$817 final_adder.U$$784/A final_adder.U$$737/X final_adder.U$$705/X
+ VGND VGND VPWR VPWR final_adder.U$$817/X sky130_fd_sc_hd__a21o_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$839 final_adder.U$$742/X final_adder.U$$807/X final_adder.U$$743/X
+ VGND VGND VPWR VPWR final_adder.U$$839/X sky130_fd_sc_hd__a21o_2
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_90_0_1928 VGND VGND VPWR VPWR dadda_fa_1_90_0/A dadda_fa_1_90_0_1928/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_165_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_95_1 dadda_fa_4_95_1/A dadda_fa_4_95_1/B dadda_fa_4_95_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_96_0/B dadda_fa_5_95_1/B sky130_fd_sc_hd__fa_1
XFILLER_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_72_0 dadda_fa_7_72_0/A dadda_fa_7_72_0/B dadda_fa_7_72_0/CIN VGND VGND
+ VPWR VPWR _369_/D _240_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_88_0 dadda_fa_4_88_0/A dadda_fa_4_88_0/B dadda_fa_4_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_89_0/A dadda_fa_5_88_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_109_3 U$$4348/X U$$4481/X input139/X VGND VGND VPWR VPWR dadda_fa_4_110_1/B
+ dadda_fa_4_109_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput370 output370/A VGND VGND VPWR VPWR o[87] sky130_fd_sc_hd__buf_2
Xoutput381 output381/A VGND VGND VPWR VPWR o[97] sky130_fd_sc_hd__buf_2
Xfanout1006 fanout1011/X VGND VGND VPWR VPWR U$$2814/A1 sky130_fd_sc_hd__buf_4
XFILLER_105_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1017 U$$4182/A1 VGND VGND VPWR VPWR U$$4043/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1028 input9/X VGND VGND VPWR VPWR U$$1221/B sky130_fd_sc_hd__buf_8
XFILLER_102_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1039 U$$479/A1 VGND VGND VPWR VPWR U$$616/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_142_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2107 U$$50/B1 U$$2107/A2 U$$739/A1 U$$2107/B2 VGND VGND VPWR VPWR U$$2108/A sky130_fd_sc_hd__a22o_1
XFILLER_16_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2118 U$$2118/A U$$2148/B VGND VGND VPWR VPWR U$$2118/X sky130_fd_sc_hd__xor2_1
XFILLER_142_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2129 U$$3499/A1 U$$2177/A2 U$$3636/B1 U$$2177/B2 VGND VGND VPWR VPWR U$$2130/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1406 U$$447/A1 U$$1414/A2 U$$447/B1 U$$1414/B2 VGND VGND VPWR VPWR U$$1407/A sky130_fd_sc_hd__a22o_1
XFILLER_35_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1417 U$$1417/A U$$1433/B VGND VGND VPWR VPWR U$$1417/X sky130_fd_sc_hd__xor2_1
XU$$1428 U$$56/B1 U$$1460/A2 U$$469/B1 U$$1460/B2 VGND VGND VPWR VPWR U$$1429/A sky130_fd_sc_hd__a22o_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1439 U$$1439/A U$$1449/B VGND VGND VPWR VPWR U$$1439/X sky130_fd_sc_hd__xor2_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_215_ _343_/CLK _215_/D VGND VGND VPWR VPWR _215_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_90_0 dadda_fa_3_90_0/A dadda_fa_3_90_0/B dadda_fa_3_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_0/B dadda_fa_4_90_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_137_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1540 U$$545/A1 VGND VGND VPWR VPWR U$$4244/A1 sky130_fd_sc_hd__buf_4
XFILLER_66_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1551 U$$3966/B1 VGND VGND VPWR VPWR U$$4240/B1 sky130_fd_sc_hd__buf_4
Xfanout1562 U$$952/A1 VGND VGND VPWR VPWR U$$3692/A1 sky130_fd_sc_hd__buf_2
XU$$4010 U$$4010/A U$$4058/B VGND VGND VPWR VPWR U$$4010/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_52_5 dadda_fa_2_52_5/A dadda_fa_2_52_5/B dadda_fa_2_52_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_2/A dadda_fa_4_52_0/A sky130_fd_sc_hd__fa_2
Xfanout1573 input121/X VGND VGND VPWR VPWR U$$950/A1 sky130_fd_sc_hd__buf_4
XU$$4021 U$$4158/A1 U$$4045/A2 U$$4295/B1 U$$4045/B2 VGND VGND VPWR VPWR U$$4022/A
+ sky130_fd_sc_hd__a22o_1
XU$$4032 U$$4032/A U$$4040/B VGND VGND VPWR VPWR U$$4032/X sky130_fd_sc_hd__xor2_1
Xfanout1584 U$$99/B VGND VGND VPWR VPWR U$$3/A sky130_fd_sc_hd__clkbuf_4
Xfanout1595 U$$2729/A1 VGND VGND VPWR VPWR U$$948/A1 sky130_fd_sc_hd__buf_4
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4043 U$$4043/A1 U$$4043/A2 U$$4043/B1 U$$4043/B2 VGND VGND VPWR VPWR U$$4044/A
+ sky130_fd_sc_hd__a22o_1
XU$$4054 U$$4054/A U$$4058/B VGND VGND VPWR VPWR U$$4054/X sky130_fd_sc_hd__xor2_1
XFILLER_19_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_45_4 dadda_fa_2_45_4/A dadda_fa_2_45_4/B dadda_fa_2_45_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_46_1/CIN dadda_fa_3_45_3/CIN sky130_fd_sc_hd__fa_1
XU$$3320 U$$989/B1 U$$3338/A2 U$$856/A1 U$$3338/B2 VGND VGND VPWR VPWR U$$3321/A sky130_fd_sc_hd__a22o_1
XU$$4065 U$$4476/A1 U$$4081/A2 U$$4478/A1 U$$4081/B2 VGND VGND VPWR VPWR U$$4066/A
+ sky130_fd_sc_hd__a22o_1
XU$$3331 U$$3331/A U$$3335/B VGND VGND VPWR VPWR U$$3331/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4076 U$$4076/A U$$4082/B VGND VGND VPWR VPWR U$$4076/X sky130_fd_sc_hd__xor2_1
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3342 U$$876/A1 U$$3390/A2 U$$878/A1 U$$3390/B2 VGND VGND VPWR VPWR U$$3343/A sky130_fd_sc_hd__a22o_1
XU$$4087 U$$4361/A1 U$$4107/A2 U$$4363/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4088/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3353 U$$3353/A U$$3424/A VGND VGND VPWR VPWR U$$3353/X sky130_fd_sc_hd__xor2_1
XU$$4098 U$$4098/A U$$4098/B VGND VGND VPWR VPWR U$$4098/X sky130_fd_sc_hd__xor2_1
XU$$3364 U$$3636/B1 U$$3372/A2 U$$3638/B1 U$$3372/B2 VGND VGND VPWR VPWR U$$3365/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_38_3 U$$2344/X U$$2477/X U$$2610/X VGND VGND VPWR VPWR dadda_fa_3_39_1/B
+ dadda_fa_3_38_3/B sky130_fd_sc_hd__fa_1
XFILLER_34_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2630 U$$2630/A U$$2668/B VGND VGND VPWR VPWR U$$2630/X sky130_fd_sc_hd__xor2_1
XU$$3375 U$$3375/A U$$3425/A VGND VGND VPWR VPWR U$$3375/X sky130_fd_sc_hd__xor2_1
XU$$3386 U$$4345/A1 U$$3416/A2 U$$4482/B1 U$$3416/B2 VGND VGND VPWR VPWR U$$3387/A
+ sky130_fd_sc_hd__a22o_1
XU$$2641 U$$4011/A1 U$$2679/A2 U$$2780/A1 U$$2679/B2 VGND VGND VPWR VPWR U$$2642/A
+ sky130_fd_sc_hd__a22o_1
XU$$3397 U$$3397/A U$$3417/B VGND VGND VPWR VPWR U$$3397/X sky130_fd_sc_hd__xor2_1
XU$$2652 U$$2652/A U$$2668/B VGND VGND VPWR VPWR U$$2652/X sky130_fd_sc_hd__xor2_1
XU$$2663 U$$4442/B1 U$$2707/A2 U$$4309/A1 U$$2707/B2 VGND VGND VPWR VPWR U$$2664/A
+ sky130_fd_sc_hd__a22o_1
XU$$2674 U$$2674/A U$$2740/A VGND VGND VPWR VPWR U$$2674/X sky130_fd_sc_hd__xor2_1
XU$$1940 U$$979/B1 U$$1980/A2 U$$3447/B1 U$$1980/B2 VGND VGND VPWR VPWR U$$1941/A
+ sky130_fd_sc_hd__a22o_1
XU$$2685 U$$4464/B1 U$$2737/A2 U$$4331/A1 U$$2737/B2 VGND VGND VPWR VPWR U$$2686/A
+ sky130_fd_sc_hd__a22o_1
XU$$1951 U$$1951/A U$$2007/B VGND VGND VPWR VPWR U$$1951/X sky130_fd_sc_hd__xor2_1
XU$$2696 U$$2696/A U$$2708/B VGND VGND VPWR VPWR U$$2696/X sky130_fd_sc_hd__xor2_1
XFILLER_61_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1962 U$$3056/B1 U$$1964/A2 U$$2923/A1 U$$1964/B2 VGND VGND VPWR VPWR U$$1963/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1973 U$$1973/A U$$1981/B VGND VGND VPWR VPWR U$$1973/X sky130_fd_sc_hd__xor2_1
XU$$1984 U$$612/B1 U$$2014/A2 U$$479/A1 U$$2014/B2 VGND VGND VPWR VPWR U$$1985/A sky130_fd_sc_hd__a22o_1
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1995 U$$1995/A U$$2031/B VGND VGND VPWR VPWR U$$1995/X sky130_fd_sc_hd__xor2_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput109 b[4] VGND VGND VPWR VPWR input109/X sky130_fd_sc_hd__buf_4
XFILLER_130_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$603 final_adder.U$$602/B final_adder.U$$487/X final_adder.U$$479/X
+ VGND VGND VPWR VPWR final_adder.U$$603/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$614 final_adder.U$$614/A final_adder.U$$614/B VGND VGND VPWR VPWR
+ final_adder.U$$718/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$625 final_adder.U$$616/A final_adder.U$$255/X final_adder.U$$501/X
+ VGND VGND VPWR VPWR final_adder.U$$625/X sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$636 final_adder.U$$652/B final_adder.U$$636/B VGND VGND VPWR VPWR
+ final_adder.U$$748/B sky130_fd_sc_hd__and2_1
XFILLER_99_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$647 final_adder.U$$646/B final_adder.U$$543/X final_adder.U$$527/X
+ VGND VGND VPWR VPWR final_adder.U$$647/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$658 final_adder.U$$674/B final_adder.U$$658/B VGND VGND VPWR VPWR
+ final_adder.U$$770/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$669 final_adder.U$$668/B final_adder.U$$565/X final_adder.U$$549/X
+ VGND VGND VPWR VPWR final_adder.U$$669/X sky130_fd_sc_hd__a21o_1
XU$$508 U$$508/A U$$522/B VGND VGND VPWR VPWR U$$508/X sky130_fd_sc_hd__xor2_1
XU$$519 U$$654/B1 U$$545/A2 U$$521/A1 U$$545/B2 VGND VGND VPWR VPWR U$$520/A sky130_fd_sc_hd__a22o_1
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$80 U$$80/A1 U$$80/A2 U$$80/B1 U$$80/B2 VGND VGND VPWR VPWR U$$81/A sky130_fd_sc_hd__a22o_1
XU$$91 U$$91/A U$$97/B VGND VGND VPWR VPWR U$$91/X sky130_fd_sc_hd__xor2_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4423_1859 VGND VGND VPWR VPWR U$$4423_1859/HI U$$4423/B sky130_fd_sc_hd__conb_1
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_107_0 U$$3413/X U$$3546/X U$$3679/X VGND VGND VPWR VPWR dadda_fa_4_108_0/B
+ dadda_fa_4_107_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_55_3 dadda_fa_3_55_3/A dadda_fa_3_55_3/B dadda_fa_3_55_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_1/B dadda_fa_4_55_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_102_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_48_2 dadda_fa_3_48_2/A dadda_fa_3_48_2/B dadda_fa_3_48_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_1/A dadda_fa_4_48_2/B sky130_fd_sc_hd__fa_1
XFILLER_46_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_18_0 dadda_fa_6_18_0/A dadda_fa_6_18_0/B dadda_fa_6_18_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_19_0/B dadda_fa_7_18_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_62_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1203 U$$1203/A U$$1233/A VGND VGND VPWR VPWR U$$1203/X sky130_fd_sc_hd__xor2_1
XFILLER_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1214 U$$253/B1 U$$1218/A2 U$$120/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1215/A sky130_fd_sc_hd__a22o_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1225 U$$1225/A U$$1227/B VGND VGND VPWR VPWR U$$1225/X sky130_fd_sc_hd__xor2_1
XU$$1236 U$$1370/A U$$1236/B VGND VGND VPWR VPWR U$$1236/X sky130_fd_sc_hd__and2_1
XU$$1247 U$$2480/A1 U$$1311/A2 U$$3030/A1 U$$1311/B2 VGND VGND VPWR VPWR U$$1248/A
+ sky130_fd_sc_hd__a22o_1
XU$$1258 U$$1258/A U$$1294/B VGND VGND VPWR VPWR U$$1258/X sky130_fd_sc_hd__xor2_1
XFILLER_71_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1269 U$$36/A1 U$$1311/A2 U$$38/A1 U$$1311/B2 VGND VGND VPWR VPWR U$$1270/A sky130_fd_sc_hd__a22o_1
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1030 final_adder.U$$6/SUM final_adder.U$$505/X VGND VGND VPWR VPWR
+ output351/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1041 final_adder.U$$238/B final_adder.U$$1041/B VGND VGND VPWR VPWR
+ output293/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1052 final_adder.U$$226/A final_adder.U$$727/X VGND VGND VPWR VPWR
+ output305/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1063 final_adder.U$$216/B final_adder.U$$987/X VGND VGND VPWR VPWR
+ output317/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1074 final_adder.U$$204/A final_adder.U$$817/X VGND VGND VPWR VPWR
+ output330/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1085 final_adder.U$$194/B final_adder.U$$965/X VGND VGND VPWR VPWR
+ output342/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1096 final_adder.U$$182/A final_adder.U$$891/X VGND VGND VPWR VPWR
+ output354/A sky130_fd_sc_hd__xor2_1
XFILLER_171_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_50_2 dadda_fa_2_50_2/A dadda_fa_2_50_2/B dadda_fa_2_50_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_1/A dadda_fa_3_50_3/A sky130_fd_sc_hd__fa_1
XFILLER_78_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1370 U$$3119/B VGND VGND VPWR VPWR U$$3150/A sky130_fd_sc_hd__buf_6
Xfanout1381 U$$2990/B VGND VGND VPWR VPWR U$$2986/B sky130_fd_sc_hd__buf_6
Xfanout1392 U$$260/B VGND VGND VPWR VPWR U$$230/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_43_1 U$$2354/X U$$2487/X U$$2620/X VGND VGND VPWR VPWR dadda_fa_3_44_0/CIN
+ dadda_fa_3_43_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_20_0 dadda_fa_5_20_0/A dadda_fa_5_20_0/B dadda_fa_5_20_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_21_0/A dadda_fa_6_20_0/CIN sky130_fd_sc_hd__fa_1
XU$$3150 U$$3150/A VGND VGND VPWR VPWR U$$3150/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_2_36_0 U$$744/X U$$877/X U$$1010/X VGND VGND VPWR VPWR dadda_fa_3_37_0/B
+ dadda_fa_3_36_2/B sky130_fd_sc_hd__fa_1
XU$$3161 U$$3296/B1 U$$3199/A2 U$$3163/A1 U$$3199/B2 VGND VGND VPWR VPWR U$$3162/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3172 U$$3172/A U$$3210/B VGND VGND VPWR VPWR U$$3172/X sky130_fd_sc_hd__xor2_1
XFILLER_53_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3183 U$$852/B1 U$$3207/A2 U$$854/B1 U$$3207/B2 VGND VGND VPWR VPWR U$$3184/A sky130_fd_sc_hd__a22o_1
XU$$3194 U$$3194/A U$$3196/B VGND VGND VPWR VPWR U$$3194/X sky130_fd_sc_hd__xor2_1
XU$$2460 U$$2460/A U$$2465/A VGND VGND VPWR VPWR U$$2460/X sky130_fd_sc_hd__xor2_1
XU$$2471 U$$2469/B U$$2466/A input30/X U$$2466/Y VGND VGND VPWR VPWR U$$2471/X sky130_fd_sc_hd__a22o_1
XFILLER_146_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2482 U$$3850/B1 U$$2540/A2 U$$4402/A1 U$$2540/B2 VGND VGND VPWR VPWR U$$2483/A
+ sky130_fd_sc_hd__a22o_1
XU$$2493 U$$2493/A U$$2529/B VGND VGND VPWR VPWR U$$2493/X sky130_fd_sc_hd__xor2_1
XU$$1770 U$$2179/B1 U$$1774/A2 U$$2183/A1 U$$1774/B2 VGND VGND VPWR VPWR U$$1771/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1781 U$$1781/A VGND VGND VPWR VPWR U$$1781/Y sky130_fd_sc_hd__inv_1
XU$$1792 U$$1792/A U$$1828/B VGND VGND VPWR VPWR U$$1792/X sky130_fd_sc_hd__xor2_1
Xinput80 b[23] VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__buf_4
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput91 b[33] VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_88_3 U$$2843/X U$$2976/X U$$3109/X VGND VGND VPWR VPWR dadda_fa_2_89_4/B
+ dadda_fa_2_88_5/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_4_65_2 dadda_fa_4_65_2/A dadda_fa_4_65_2/B dadda_fa_4_65_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_66_0/CIN dadda_fa_5_65_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_153_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_58_1 dadda_fa_4_58_1/A dadda_fa_4_58_1/B dadda_fa_4_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_59_0/B dadda_fa_5_58_1/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$400 final_adder.U$$404/B final_adder.U$$400/B VGND VGND VPWR VPWR
+ final_adder.U$$524/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$411 final_adder.U$$410/B final_adder.U$$289/X final_adder.U$$285/X
+ VGND VGND VPWR VPWR final_adder.U$$411/X sky130_fd_sc_hd__a21o_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_35_0 dadda_fa_7_35_0/A dadda_fa_7_35_0/B dadda_fa_7_35_0/CIN VGND VGND
+ VPWR VPWR _332_/D _203_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$422 final_adder.U$$426/B final_adder.U$$422/B VGND VGND VPWR VPWR
+ final_adder.U$$546/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$433 final_adder.U$$432/B final_adder.U$$311/X final_adder.U$$307/X
+ VGND VGND VPWR VPWR final_adder.U$$433/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$444 final_adder.U$$448/B final_adder.U$$444/B VGND VGND VPWR VPWR
+ final_adder.U$$568/B sky130_fd_sc_hd__and2_1
XFILLER_123_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$455 final_adder.U$$454/B final_adder.U$$333/X final_adder.U$$329/X
+ VGND VGND VPWR VPWR final_adder.U$$455/X sky130_fd_sc_hd__a21o_1
XFILLER_45_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$466 final_adder.U$$470/B final_adder.U$$466/B VGND VGND VPWR VPWR
+ final_adder.U$$590/B sky130_fd_sc_hd__and2_1
XFILLER_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$305 U$$305/A U$$339/B VGND VGND VPWR VPWR U$$305/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$477 final_adder.U$$476/B final_adder.U$$355/X final_adder.U$$351/X
+ VGND VGND VPWR VPWR final_adder.U$$477/X sky130_fd_sc_hd__a21o_1
XU$$316 U$$40/B1 U$$338/A2 U$$316/B1 U$$338/B2 VGND VGND VPWR VPWR U$$317/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$488 final_adder.U$$492/B final_adder.U$$488/B VGND VGND VPWR VPWR
+ final_adder.U$$612/B sky130_fd_sc_hd__and2_1
XU$$327 U$$327/A U$$363/B VGND VGND VPWR VPWR U$$327/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$499 final_adder.U$$498/B final_adder.U$$377/X final_adder.U$$373/X
+ VGND VGND VPWR VPWR final_adder.U$$499/X sky130_fd_sc_hd__a21o_1
XU$$338 U$$747/B1 U$$338/A2 U$$749/B1 U$$338/B2 VGND VGND VPWR VPWR U$$339/A sky130_fd_sc_hd__a22o_1
XU$$349 U$$349/A U$$353/B VGND VGND VPWR VPWR U$$349/X sky130_fd_sc_hd__xor2_1
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_60_1 dadda_fa_3_60_1/A dadda_fa_3_60_1/B dadda_fa_3_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_0/CIN dadda_fa_4_60_2/A sky130_fd_sc_hd__fa_1
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_53_0 dadda_fa_3_53_0/A dadda_fa_3_53_0/B dadda_fa_3_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_0/B dadda_fa_4_53_1/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_0_69_0 U$$410/Y U$$544/X U$$677/X VGND VGND VPWR VPWR dadda_fa_1_70_6/A
+ dadda_fa_1_69_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$850 U$$850/A1 U$$898/A2 U$$989/A1 U$$898/B2 VGND VGND VPWR VPWR U$$851/A sky130_fd_sc_hd__a22o_1
XU$$861 U$$861/A U$$895/B VGND VGND VPWR VPWR U$$861/X sky130_fd_sc_hd__xor2_1
XU$$1000 U$$999/X U$$1062/B VGND VGND VPWR VPWR U$$1000/X sky130_fd_sc_hd__xor2_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1011 U$$50/B1 U$$979/A2 U$$739/A1 U$$979/B2 VGND VGND VPWR VPWR U$$1012/A sky130_fd_sc_hd__a22o_1
XU$$872 U$$872/A1 U$$876/A2 U$$874/A1 U$$876/B2 VGND VGND VPWR VPWR U$$873/A sky130_fd_sc_hd__a22o_1
XU$$1022 U$$1022/A U$$998/B VGND VGND VPWR VPWR U$$1022/X sky130_fd_sc_hd__xor2_1
XU$$883 U$$883/A U$$907/B VGND VGND VPWR VPWR U$$883/X sky130_fd_sc_hd__xor2_1
XU$$894 U$$894/A1 U$$898/A2 U$$896/A1 U$$898/B2 VGND VGND VPWR VPWR U$$895/A sky130_fd_sc_hd__a22o_1
XU$$1033 U$$896/A1 U$$1075/A2 U$$898/A1 U$$1075/B2 VGND VGND VPWR VPWR U$$1034/A sky130_fd_sc_hd__a22o_1
XU$$4445_1870 VGND VGND VPWR VPWR U$$4445_1870/HI U$$4445/B sky130_fd_sc_hd__conb_1
XU$$1044 U$$1044/A U$$1046/B VGND VGND VPWR VPWR U$$1044/X sky130_fd_sc_hd__xor2_1
XU$$1055 U$$96/A1 U$$1075/A2 U$$98/A1 U$$1075/B2 VGND VGND VPWR VPWR U$$1056/A sky130_fd_sc_hd__a22o_1
XU$$1066 U$$1066/A U$$962/A VGND VGND VPWR VPWR U$$1066/X sky130_fd_sc_hd__xor2_1
XU$$1077 U$$803/A1 U$$1093/A2 U$$805/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1078/A sky130_fd_sc_hd__a22o_1
XFILLER_32_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1088 U$$1088/A U$$1088/B VGND VGND VPWR VPWR U$$1088/X sky130_fd_sc_hd__xor2_1
XU$$1099 U$$1233/A U$$1099/B VGND VGND VPWR VPWR U$$1099/X sky130_fd_sc_hd__and2_1
XFILLER_31_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_110_0 dadda_fa_7_110_0/A dadda_fa_7_110_0/B dadda_fa_7_110_0/CIN VGND
+ VGND VPWR VPWR _407_/D _278_/D sky130_fd_sc_hd__fa_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_98_2 U$$3129/X U$$3262/X U$$3395/X VGND VGND VPWR VPWR dadda_fa_3_99_1/B
+ dadda_fa_3_98_3/A sky130_fd_sc_hd__fa_1
XFILLER_160_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_75_1 dadda_fa_5_75_1/A dadda_fa_5_75_1/B dadda_fa_5_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_76_0/B dadda_fa_7_75_0/A sky130_fd_sc_hd__fa_1
XFILLER_137_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_68_0 dadda_fa_5_68_0/A dadda_fa_5_68_0/B dadda_fa_5_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_69_0/A dadda_fa_6_68_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_98_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout607 U$$1760/A2 VGND VGND VPWR VPWR U$$1720/A2 sky130_fd_sc_hd__buf_4
Xfanout618 U$$1625/A2 VGND VGND VPWR VPWR U$$1635/A2 sky130_fd_sc_hd__clkbuf_4
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout629 U$$1460/A2 VGND VGND VPWR VPWR U$$1426/A2 sky130_fd_sc_hd__buf_4
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_8 dadda_fa_1_67_8/A dadda_fa_1_67_8/B dadda_fa_1_67_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_68_3/A dadda_fa_3_67_0/A sky130_fd_sc_hd__fa_1
XFILLER_101_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_7_0 dadda_fa_6_7_0/A dadda_fa_6_7_0/B dadda_fa_6_7_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_8_0/B dadda_fa_7_7_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_23_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2290 U$$3249/A1 U$$2326/A2 U$$3249/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2291/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_93_1 U$$2454/X U$$2587/X U$$2720/X VGND VGND VPWR VPWR dadda_fa_2_94_5/B
+ dadda_fa_3_93_0/A sky130_fd_sc_hd__fa_1
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_70_0 dadda_fa_4_70_0/A dadda_fa_4_70_0/B dadda_fa_4_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_71_0/A dadda_fa_5_70_1/A sky130_fd_sc_hd__fa_1
XFILLER_104_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_86_0 dadda_fa_1_86_0/A U$$1642/X U$$1775/X VGND VGND VPWR VPWR dadda_fa_2_87_2/CIN
+ dadda_fa_2_86_4/B sky130_fd_sc_hd__fa_1
XFILLER_49_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_2_106_1 U$$3278/X U$$3411/X VGND VGND VPWR VPWR dadda_fa_3_107_3/CIN dadda_fa_4_106_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_40_1003 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$230 final_adder.U$$230/A final_adder.U$$230/B VGND VGND VPWR VPWR
+ final_adder.U$$358/B sky130_fd_sc_hd__and2_1
XU$$3908 U$$4043/B1 U$$3912/A2 U$$3908/B1 U$$3912/B2 VGND VGND VPWR VPWR U$$3909/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$241 final_adder.U$$240/B final_adder.U$$241/A2 final_adder.U$$241/B1
+ VGND VGND VPWR VPWR final_adder.U$$241/X sky130_fd_sc_hd__a21o_1
XU$$3919 U$$3919/A U$$3949/B VGND VGND VPWR VPWR U$$3919/X sky130_fd_sc_hd__xor2_1
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$252 final_adder.U$$252/A final_adder.U$$3/SUM VGND VGND VPWR VPWR
+ final_adder.U$$378/A sky130_fd_sc_hd__and2_1
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$263 final_adder.U$$262/B final_adder.U$$137/X final_adder.U$$135/X
+ VGND VGND VPWR VPWR final_adder.U$$263/X sky130_fd_sc_hd__a21o_1
XFILLER_18_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$102 U$$924/A1 U$$102/A2 U$$926/A1 U$$102/B2 VGND VGND VPWR VPWR U$$103/A sky130_fd_sc_hd__a22o_1
XFILLER_100_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$274 final_adder.U$$276/B final_adder.U$$274/B VGND VGND VPWR VPWR
+ final_adder.U$$400/B sky130_fd_sc_hd__and2_1
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$113 U$$113/A U$$121/B VGND VGND VPWR VPWR U$$113/X sky130_fd_sc_hd__xor2_1
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$285 final_adder.U$$284/B final_adder.U$$159/X final_adder.U$$157/X
+ VGND VGND VPWR VPWR final_adder.U$$285/X sky130_fd_sc_hd__a21o_1
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$124 U$$672/A1 U$$98/A2 U$$672/B1 U$$98/B2 VGND VGND VPWR VPWR U$$125/A sky130_fd_sc_hd__a22o_1
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$296 final_adder.U$$298/B final_adder.U$$296/B VGND VGND VPWR VPWR
+ final_adder.U$$422/B sky130_fd_sc_hd__and2_1
XU$$135 U$$135/A U$$3/A VGND VGND VPWR VPWR U$$135/X sky130_fd_sc_hd__xor2_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$146 U$$146/A U$$180/B VGND VGND VPWR VPWR U$$146/X sky130_fd_sc_hd__xor2_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$157 U$$20/A1 U$$179/A2 U$$22/A1 U$$179/B2 VGND VGND VPWR VPWR U$$158/A sky130_fd_sc_hd__a22o_1
XU$$168 U$$168/A U$$210/B VGND VGND VPWR VPWR U$$168/X sky130_fd_sc_hd__xor2_1
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$179 U$$42/A1 U$$179/A2 U$$44/A1 U$$179/B2 VGND VGND VPWR VPWR U$$180/A sky130_fd_sc_hd__a22o_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_394_ _397_/CLK _394_/D VGND VGND VPWR VPWR _394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_85_0 dadda_fa_6_85_0/A dadda_fa_6_85_0/B dadda_fa_6_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_86_0/B dadda_fa_7_85_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4475_1885 VGND VGND VPWR VPWR U$$4475_1885/HI U$$4475/B sky130_fd_sc_hd__conb_1
XFILLER_5_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$680 U$$954/A1 U$$682/A2 U$$956/A1 U$$682/B2 VGND VGND VPWR VPWR U$$681/A sky130_fd_sc_hd__a22o_1
XU$$691 U$$691/A1 U$$743/A2 U$$965/B1 U$$743/B2 VGND VGND VPWR VPWR U$$692/A sky130_fd_sc_hd__a22o_1
XFILLER_17_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_919 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout404 U$$771/A2 VGND VGND VPWR VPWR U$$743/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_160_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout415 U$$552/X VGND VGND VPWR VPWR U$$642/A2 sky130_fd_sc_hd__buf_4
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout426 U$$543/A2 VGND VGND VPWR VPWR U$$501/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_72_6 U$$4407/X input226/X dadda_fa_1_72_6/CIN VGND VGND VPWR VPWR dadda_fa_2_73_2/B
+ dadda_fa_2_72_5/B sky130_fd_sc_hd__fa_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout437 U$$4114/X VGND VGND VPWR VPWR U$$4236/A2 sky130_fd_sc_hd__clkbuf_2
Xfanout448 U$$102/A2 VGND VGND VPWR VPWR U$$120/A2 sky130_fd_sc_hd__buf_6
XFILLER_113_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout459 U$$3872/A2 VGND VGND VPWR VPWR U$$3892/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_65_5 input218/X dadda_fa_1_65_5/B dadda_fa_1_65_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_66_2/A dadda_fa_2_65_5/A sky130_fd_sc_hd__fa_1
XFILLER_86_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_58_4 U$$3182/X U$$3315/X U$$3448/X VGND VGND VPWR VPWR dadda_fa_2_59_1/CIN
+ dadda_fa_2_58_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_28_2 dadda_fa_4_28_2/A dadda_fa_4_28_2/B dadda_fa_4_28_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_29_0/CIN dadda_fa_5_28_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_918 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout960 U$$3509/A1 VGND VGND VPWR VPWR U$$3370/B1 sky130_fd_sc_hd__buf_4
XU$$4406 U$$4406/A1 U$$4388/X U$$4408/A1 U$$4458/B2 VGND VGND VPWR VPWR U$$4407/A
+ sky130_fd_sc_hd__a22o_1
XU$$4417 U$$4417/A U$$4417/B VGND VGND VPWR VPWR U$$4417/X sky130_fd_sc_hd__xor2_1
Xfanout971 fanout975/X VGND VGND VPWR VPWR U$$82/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_38_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4428 U$$4428/A1 U$$4388/X U$$4430/A1 U$$4428/B2 VGND VGND VPWR VPWR U$$4429/A
+ sky130_fd_sc_hd__a22o_1
Xfanout982 fanout984/X VGND VGND VPWR VPWR U$$3916/A1 sky130_fd_sc_hd__buf_6
Xfanout993 input93/X VGND VGND VPWR VPWR fanout993/X sky130_fd_sc_hd__buf_8
XU$$4439 U$$4439/A U$$4439/B VGND VGND VPWR VPWR U$$4439/X sky130_fd_sc_hd__xor2_1
XU$$3705 U$$3705/A1 U$$3791/A2 U$$3979/B1 U$$3791/B2 VGND VGND VPWR VPWR U$$3706/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3716 U$$3716/A U$$3740/B VGND VGND VPWR VPWR U$$3716/X sky130_fd_sc_hd__xor2_1
XU$$3727 U$$3999/B1 U$$3757/A2 U$$4001/B1 U$$3757/B2 VGND VGND VPWR VPWR U$$3728/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3738 U$$3738/A U$$3740/B VGND VGND VPWR VPWR U$$3738/X sky130_fd_sc_hd__xor2_1
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3749 U$$4434/A1 U$$3829/A2 U$$3751/A1 U$$3829/B2 VGND VGND VPWR VPWR U$$3750/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_2 dadda_fa_3_30_2/A dadda_fa_3_30_2/B dadda_fa_3_30_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_31_1/A dadda_fa_4_30_2/B sky130_fd_sc_hd__fa_1
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_23_1 U$$718/X U$$851/X U$$984/X VGND VGND VPWR VPWR dadda_fa_4_24_0/CIN
+ dadda_fa_4_23_2/A sky130_fd_sc_hd__fa_2
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_16_0 U$$39/X U$$172/X U$$305/X VGND VGND VPWR VPWR dadda_fa_4_17_1/CIN
+ dadda_fa_4_16_2/B sky130_fd_sc_hd__fa_1
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_377_ _377_/CLK _377_/D VGND VGND VPWR VPWR _377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$691_1912 VGND VGND VPWR VPWR U$$691_1912/HI U$$691/A1 sky130_fd_sc_hd__conb_1
XFILLER_173_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_82_5 dadda_fa_2_82_5/A dadda_fa_2_82_5/B dadda_fa_2_82_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_2/A dadda_fa_4_82_0/A sky130_fd_sc_hd__fa_2
XFILLER_142_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_75_4 dadda_fa_2_75_4/A dadda_fa_2_75_4/B dadda_fa_2_75_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_1/CIN dadda_fa_3_75_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_68_3 dadda_fa_2_68_3/A dadda_fa_2_68_3/B dadda_fa_2_68_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_1/B dadda_fa_3_68_3/B sky130_fd_sc_hd__fa_1
XFILLER_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_38_1 dadda_fa_5_38_1/A dadda_fa_5_38_1/B dadda_fa_5_38_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_39_0/B dadda_fa_7_38_0/A sky130_fd_sc_hd__fa_1
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_112_1 dadda_fa_5_112_1/A dadda_fa_5_112_1/B dadda_fa_5_112_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_113_0/B dadda_fa_7_112_0/A sky130_fd_sc_hd__fa_1
XFILLER_30_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_105_0 dadda_fa_5_105_0/A dadda_fa_5_105_0/B dadda_fa_5_105_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_106_0/A dadda_fa_6_105_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_133_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_70_3 U$$3472/X U$$3605/X U$$3738/X VGND VGND VPWR VPWR dadda_fa_2_71_1/B
+ dadda_fa_2_70_4/B sky130_fd_sc_hd__fa_1
XFILLER_101_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_63_2 U$$3192/X U$$3325/X U$$3458/X VGND VGND VPWR VPWR dadda_fa_2_64_1/A
+ dadda_fa_2_63_4/A sky130_fd_sc_hd__fa_1
XFILLER_59_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_40_1 dadda_fa_4_40_1/A dadda_fa_4_40_1/B dadda_fa_4_40_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_41_0/B dadda_fa_5_40_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_56_1 U$$1582/X U$$1715/X U$$1848/X VGND VGND VPWR VPWR dadda_fa_2_57_0/CIN
+ dadda_fa_2_56_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_4_33_0 dadda_fa_4_33_0/A dadda_fa_4_33_0/B dadda_fa_4_33_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_34_0/A dadda_fa_5_33_1/A sky130_fd_sc_hd__fa_1
XFILLER_55_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_49_0 U$$105/X U$$238/X U$$371/X VGND VGND VPWR VPWR dadda_fa_2_50_0/CIN
+ dadda_fa_2_49_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_300_ _319_/CLK _300_/D VGND VGND VPWR VPWR _300_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_231_ _360_/CLK _231_/D VGND VGND VPWR VPWR _231_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_85_3 dadda_fa_3_85_3/A dadda_fa_3_85_3/B dadda_fa_3_85_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_1/B dadda_fa_4_85_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_78_2 dadda_fa_3_78_2/A dadda_fa_3_78_2/B dadda_fa_3_78_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_1/A dadda_fa_4_78_2/B sky130_fd_sc_hd__fa_1
Xfanout1700 input109/X VGND VGND VPWR VPWR U$$3713/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1711 U$$2979/B1 VGND VGND VPWR VPWR U$$2707/A1 sky130_fd_sc_hd__buf_4
XFILLER_2_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1722 input106/X VGND VGND VPWR VPWR U$$787/A1 sky130_fd_sc_hd__buf_6
Xfanout1733 U$$3249/B1 VGND VGND VPWR VPWR U$$4484/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_48_0 dadda_fa_6_48_0/A dadda_fa_6_48_0/B dadda_fa_6_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_49_0/B dadda_fa_7_48_0/CIN sky130_fd_sc_hd__fa_1
Xfanout1744 U$$505/B1 VGND VGND VPWR VPWR U$$96/A1 sky130_fd_sc_hd__buf_4
Xfanout1755 U$$3243/B1 VGND VGND VPWR VPWR U$$3106/B1 sky130_fd_sc_hd__buf_4
XFILLER_77_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4203 U$$4203/A U$$4215/B VGND VGND VPWR VPWR U$$4203/X sky130_fd_sc_hd__xor2_1
XFILLER_172_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4214 U$$4349/B1 U$$4224/A2 U$$4214/B1 U$$4224/B2 VGND VGND VPWR VPWR U$$4215/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1766 U$$914/A1 VGND VGND VPWR VPWR U$$640/A1 sky130_fd_sc_hd__buf_6
XU$$4225 U$$4225/A U$$4227/B VGND VGND VPWR VPWR U$$4225/X sky130_fd_sc_hd__xor2_1
Xfanout1777 U$$3650/B1 VGND VGND VPWR VPWR U$$4474/A1 sky130_fd_sc_hd__clkbuf_2
Xfanout790 U$$279/X VGND VGND VPWR VPWR U$$408/B2 sky130_fd_sc_hd__buf_4
XU$$4236 U$$4508/B1 U$$4236/A2 U$$4375/A1 U$$4236/B2 VGND VGND VPWR VPWR U$$4237/A
+ sky130_fd_sc_hd__a22o_1
XU$$3502 U$$3502/A U$$3506/B VGND VGND VPWR VPWR U$$3502/X sky130_fd_sc_hd__xor2_1
XU$$4247 U$$4247/A VGND VGND VPWR VPWR U$$4247/Y sky130_fd_sc_hd__inv_1
XFILLER_92_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4258 U$$4258/A U$$4292/B VGND VGND VPWR VPWR U$$4258/X sky130_fd_sc_hd__xor2_1
XFILLER_93_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3513 U$$3650/A1 U$$3557/A2 U$$3650/B1 U$$3557/B2 VGND VGND VPWR VPWR U$$3514/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4269 U$$981/A1 U$$4289/A2 U$$4271/A1 U$$4289/B2 VGND VGND VPWR VPWR U$$4270/A
+ sky130_fd_sc_hd__a22o_1
XU$$3524 U$$3524/A U$$3524/B VGND VGND VPWR VPWR U$$3524/X sky130_fd_sc_hd__xor2_1
XU$$3535 U$$4081/B1 U$$3559/A2 U$$3948/A1 U$$3559/B2 VGND VGND VPWR VPWR U$$3536/A
+ sky130_fd_sc_hd__a22o_1
XU$$2801 U$$2801/A U$$2805/B VGND VGND VPWR VPWR U$$2801/X sky130_fd_sc_hd__xor2_1
XU$$3546 U$$3546/A U$$3548/B VGND VGND VPWR VPWR U$$3546/X sky130_fd_sc_hd__xor2_1
XFILLER_18_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3557 U$$4240/B1 U$$3557/A2 U$$4107/A1 U$$3557/B2 VGND VGND VPWR VPWR U$$3558/A
+ sky130_fd_sc_hd__a22o_1
XU$$2812 U$$346/A1 U$$2812/A2 U$$2814/A1 U$$2812/B2 VGND VGND VPWR VPWR U$$2813/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2823 U$$2823/A U$$2876/A VGND VGND VPWR VPWR U$$2823/X sky130_fd_sc_hd__xor2_1
XU$$3568 U$$3568/A1 U$$3656/A2 U$$3979/B1 U$$3656/B2 VGND VGND VPWR VPWR U$$3569/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_107_2 dadda_fa_4_107_2/A dadda_fa_4_107_2/B dadda_fa_4_107_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_108_0/CIN dadda_fa_5_107_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2834 U$$3106/B1 U$$2840/A2 U$$2973/A1 U$$2840/B2 VGND VGND VPWR VPWR U$$2835/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_836 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3579 U$$3579/A U$$3615/B VGND VGND VPWR VPWR U$$3579/X sky130_fd_sc_hd__xor2_1
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2845 U$$2845/A U$$2877/A VGND VGND VPWR VPWR U$$2845/X sky130_fd_sc_hd__xor2_1
XU$$2856 U$$251/B1 U$$2856/A2 U$$2993/B1 U$$2856/B2 VGND VGND VPWR VPWR U$$2857/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2867 U$$2867/A U$$2871/B VGND VGND VPWR VPWR U$$2867/X sky130_fd_sc_hd__xor2_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2878 input37/X VGND VGND VPWR VPWR U$$2880/B sky130_fd_sc_hd__inv_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2889 U$$3163/A1 U$$2929/A2 U$$3163/B1 U$$2929/B2 VGND VGND VPWR VPWR U$$2890/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_80_2 dadda_fa_2_80_2/A dadda_fa_2_80_2/B dadda_fa_2_80_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_1/A dadda_fa_3_80_3/A sky130_fd_sc_hd__fa_1
XFILLER_69_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_73_1 dadda_fa_2_73_1/A dadda_fa_2_73_1/B dadda_fa_2_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_0/CIN dadda_fa_3_73_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_50_0 dadda_fa_5_50_0/A dadda_fa_5_50_0/B dadda_fa_5_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_51_0/A dadda_fa_6_50_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_60_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_66_0 dadda_fa_2_66_0/A dadda_fa_2_66_0/B dadda_fa_2_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_0/B dadda_fa_3_66_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$807 final_adder.U$$774/A final_adder.U$$727/X final_adder.U$$695/X
+ VGND VGND VPWR VPWR final_adder.U$$807/X sky130_fd_sc_hd__a21o_1
XFILLER_84_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$829 final_adder.U$$796/A final_adder.U$$505/X final_adder.U$$717/X
+ VGND VGND VPWR VPWR final_adder.U$$829/X sky130_fd_sc_hd__a21o_1
XFILLER_110_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 a[0] VGND VGND VPWR VPWR U$$1/A sky130_fd_sc_hd__buf_2
XFILLER_84_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_858 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_95_2 dadda_fa_4_95_2/A dadda_fa_4_95_2/B dadda_fa_4_95_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_96_0/CIN dadda_fa_5_95_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_88_1 dadda_fa_4_88_1/A dadda_fa_4_88_1/B dadda_fa_4_88_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_89_0/B dadda_fa_5_88_1/B sky130_fd_sc_hd__fa_1
XFILLER_118_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_65_0 dadda_fa_7_65_0/A dadda_fa_7_65_0/B dadda_fa_7_65_0/CIN VGND VGND
+ VPWR VPWR _362_/D _233_/D sky130_fd_sc_hd__fa_1
XFILLER_106_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput360 output360/A VGND VGND VPWR VPWR o[78] sky130_fd_sc_hd__buf_2
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput371 output371/A VGND VGND VPWR VPWR o[88] sky130_fd_sc_hd__buf_2
Xoutput382 output382/A VGND VGND VPWR VPWR o[98] sky130_fd_sc_hd__buf_2
Xfanout1007 fanout1011/X VGND VGND VPWR VPWR U$$3499/A1 sky130_fd_sc_hd__buf_6
XFILLER_59_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1018 U$$4182/A1 VGND VGND VPWR VPWR U$$4456/A1 sky130_fd_sc_hd__buf_4
Xfanout1029 U$$70/A1 VGND VGND VPWR VPWR U$$892/A1 sky130_fd_sc_hd__buf_4
XFILLER_87_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_39_clk _218_/CLK VGND VGND VPWR VPWR _360_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_142_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2108 U$$2108/A U$$2148/B VGND VGND VPWR VPWR U$$2108/X sky130_fd_sc_hd__xor2_1
XU$$2119 U$$612/A1 U$$2059/X U$$612/B1 U$$2060/X VGND VGND VPWR VPWR U$$2120/A sky130_fd_sc_hd__a22o_1
XFILLER_15_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1407 U$$1407/A U$$1415/B VGND VGND VPWR VPWR U$$1407/X sky130_fd_sc_hd__xor2_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1418 U$$868/B1 U$$1426/A2 U$$735/A1 U$$1426/B2 VGND VGND VPWR VPWR U$$1419/A sky130_fd_sc_hd__a22o_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1429 U$$1429/A U$$1461/B VGND VGND VPWR VPWR U$$1429/X sky130_fd_sc_hd__xor2_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_214_ _343_/CLK _214_/D VGND VGND VPWR VPWR _214_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_168_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_90_1 dadda_fa_3_90_1/A dadda_fa_3_90_1/B dadda_fa_3_90_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_0/CIN dadda_fa_4_90_2/A sky130_fd_sc_hd__fa_1
XFILLER_171_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_83_0 dadda_fa_3_83_0/A dadda_fa_3_83_0/B dadda_fa_3_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_0/B dadda_fa_4_83_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_125_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1530 input126/X VGND VGND VPWR VPWR U$$4406/A1 sky130_fd_sc_hd__buf_4
XFILLER_78_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1541 input124/X VGND VGND VPWR VPWR U$$545/A1 sky130_fd_sc_hd__buf_4
XU$$4000 U$$4000/A U$$4026/B VGND VGND VPWR VPWR U$$4000/X sky130_fd_sc_hd__xor2_1
Xfanout1552 U$$3692/B1 VGND VGND VPWR VPWR U$$3966/B1 sky130_fd_sc_hd__buf_2
Xfanout1563 U$$4514/A1 VGND VGND VPWR VPWR U$$952/A1 sky130_fd_sc_hd__buf_6
XFILLER_66_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4011 U$$4011/A1 U$$4057/A2 U$$4150/A1 U$$4057/B2 VGND VGND VPWR VPWR U$$4012/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1574 U$$3030/B1 VGND VGND VPWR VPWR U$$2758/A1 sky130_fd_sc_hd__clkbuf_4
XU$$4022 U$$4022/A U$$4040/B VGND VGND VPWR VPWR U$$4022/X sky130_fd_sc_hd__xor2_1
XU$$4033 U$$4307/A1 U$$4045/A2 U$$4307/B1 U$$4045/B2 VGND VGND VPWR VPWR U$$4034/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1585 U$$127/B VGND VGND VPWR VPWR U$$99/B sky130_fd_sc_hd__buf_6
XU$$4044 U$$4044/A U$$4110/A VGND VGND VPWR VPWR U$$4044/X sky130_fd_sc_hd__xor2_1
Xfanout1596 U$$4234/B1 VGND VGND VPWR VPWR U$$4508/B1 sky130_fd_sc_hd__buf_4
XFILLER_54_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4055 U$$4464/B1 U$$4057/A2 U$$4331/A1 U$$4057/B2 VGND VGND VPWR VPWR U$$4056/A
+ sky130_fd_sc_hd__a22o_1
XU$$3310 U$$4406/A1 U$$3390/A2 U$$4408/A1 U$$3390/B2 VGND VGND VPWR VPWR U$$3311/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_45_5 dadda_fa_2_45_5/A dadda_fa_2_45_5/B dadda_fa_2_45_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_46_2/A dadda_fa_4_45_0/A sky130_fd_sc_hd__fa_1
XU$$3321 U$$3321/A U$$3335/B VGND VGND VPWR VPWR U$$3321/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_112_0 U$$4354/X U$$4487/X input143/X VGND VGND VPWR VPWR dadda_fa_5_113_0/A
+ dadda_fa_5_112_1/A sky130_fd_sc_hd__fa_1
XU$$4066 U$$4066/A U$$4082/B VGND VGND VPWR VPWR U$$4066/X sky130_fd_sc_hd__xor2_1
XU$$3332 U$$4428/A1 U$$3372/A2 U$$4430/A1 U$$3372/B2 VGND VGND VPWR VPWR U$$3333/A
+ sky130_fd_sc_hd__a22o_1
XU$$4077 U$$4349/B1 U$$4081/A2 U$$4214/B1 U$$4081/B2 VGND VGND VPWR VPWR U$$4078/A
+ sky130_fd_sc_hd__a22o_1
XU$$3343 U$$3343/A U$$3349/B VGND VGND VPWR VPWR U$$3343/X sky130_fd_sc_hd__xor2_1
XU$$4088 U$$4088/A U$$4098/B VGND VGND VPWR VPWR U$$4088/X sky130_fd_sc_hd__xor2_1
XU$$3354 U$$3628/A1 U$$3378/A2 U$$3628/B1 U$$3378/B2 VGND VGND VPWR VPWR U$$3355/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_38_4 U$$2678/B input188/X dadda_fa_2_38_4/CIN VGND VGND VPWR VPWR dadda_fa_3_39_1/CIN
+ dadda_fa_3_38_3/CIN sky130_fd_sc_hd__fa_1
XU$$4099 U$$4508/B1 U$$4105/A2 U$$4375/A1 U$$4105/B2 VGND VGND VPWR VPWR U$$4100/A
+ sky130_fd_sc_hd__a22o_1
XU$$2620 U$$2620/A U$$2662/B VGND VGND VPWR VPWR U$$2620/X sky130_fd_sc_hd__xor2_1
XU$$3365 U$$3365/A U$$3373/B VGND VGND VPWR VPWR U$$3365/X sky130_fd_sc_hd__xor2_1
XU$$3376 U$$3376/A1 U$$3378/A2 U$$3376/B1 U$$3378/B2 VGND VGND VPWR VPWR U$$3377/A
+ sky130_fd_sc_hd__a22o_1
XU$$2631 U$$2631/A1 U$$2667/A2 U$$2631/B1 U$$2667/B2 VGND VGND VPWR VPWR U$$2632/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3387 U$$3387/A U$$3417/B VGND VGND VPWR VPWR U$$3387/X sky130_fd_sc_hd__xor2_1
XU$$2642 U$$2642/A U$$2724/B VGND VGND VPWR VPWR U$$2642/X sky130_fd_sc_hd__xor2_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2653 U$$3338/A1 U$$2667/A2 U$$735/B1 U$$2667/B2 VGND VGND VPWR VPWR U$$2654/A
+ sky130_fd_sc_hd__a22o_1
XU$$3398 U$$4081/B1 U$$3418/A2 U$$3948/A1 U$$3418/B2 VGND VGND VPWR VPWR U$$3399/A
+ sky130_fd_sc_hd__a22o_1
XU$$4409_1852 VGND VGND VPWR VPWR U$$4409_1852/HI U$$4409/B sky130_fd_sc_hd__conb_1
XU$$2664 U$$2664/A U$$2708/B VGND VGND VPWR VPWR U$$2664/X sky130_fd_sc_hd__xor2_1
XU$$1930 U$$2887/B1 U$$2006/A2 U$$2754/A1 U$$2006/B2 VGND VGND VPWR VPWR U$$1931/A
+ sky130_fd_sc_hd__a22o_1
XU$$2675 U$$4456/A1 U$$2733/A2 U$$4456/B1 U$$2733/B2 VGND VGND VPWR VPWR U$$2676/A
+ sky130_fd_sc_hd__a22o_1
XU$$1941 U$$1941/A U$$1981/B VGND VGND VPWR VPWR U$$1941/X sky130_fd_sc_hd__xor2_1
XU$$2686 U$$2686/A U$$2738/B VGND VGND VPWR VPWR U$$2686/X sky130_fd_sc_hd__xor2_1
XU$$1952 U$$993/A1 U$$1964/A2 U$$995/A1 U$$1964/B2 VGND VGND VPWR VPWR U$$1953/A sky130_fd_sc_hd__a22o_1
XU$$2697 U$$3106/B1 U$$2707/A2 U$$2973/A1 U$$2707/B2 VGND VGND VPWR VPWR U$$2698/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1963 U$$1963/A U$$1963/B VGND VGND VPWR VPWR U$$1963/X sky130_fd_sc_hd__xor2_1
XFILLER_61_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1974 U$$741/A1 U$$1986/A2 U$$880/A1 U$$1986/B2 VGND VGND VPWR VPWR U$$1975/A sky130_fd_sc_hd__a22o_1
XFILLER_21_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1985 U$$1985/A U$$2015/B VGND VGND VPWR VPWR U$$1985/X sky130_fd_sc_hd__xor2_1
XU$$1996 U$$3638/B1 U$$2046/A2 U$$3503/B1 U$$2046/B2 VGND VGND VPWR VPWR U$$1997/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_98_0 dadda_fa_5_98_0/A dadda_fa_5_98_0/B dadda_fa_5_98_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_99_0/A dadda_fa_6_98_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_147_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$604 final_adder.U$$612/B final_adder.U$$604/B VGND VGND VPWR VPWR
+ final_adder.U$$708/A sky130_fd_sc_hd__and2_1
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$615 final_adder.U$$614/B final_adder.U$$499/X final_adder.U$$491/X
+ VGND VGND VPWR VPWR final_adder.U$$615/X sky130_fd_sc_hd__a21o_1
XFILLER_69_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$637 final_adder.U$$636/B final_adder.U$$533/X final_adder.U$$517/X
+ VGND VGND VPWR VPWR final_adder.U$$637/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$648 final_adder.U$$664/B final_adder.U$$648/B VGND VGND VPWR VPWR
+ final_adder.U$$760/B sky130_fd_sc_hd__and2_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$659 final_adder.U$$658/B final_adder.U$$555/X final_adder.U$$539/X
+ VGND VGND VPWR VPWR final_adder.U$$659/X sky130_fd_sc_hd__a21o_1
XFILLER_45_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$509 U$$783/A1 U$$545/A2 U$$783/B1 U$$545/B2 VGND VGND VPWR VPWR U$$510/A sky130_fd_sc_hd__a22o_1
XFILLER_65_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$70 U$$70/A1 U$$86/A2 U$$70/B1 U$$86/B2 VGND VGND VPWR VPWR U$$71/A sky130_fd_sc_hd__a22o_1
XFILLER_25_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$81 U$$81/A U$$81/B VGND VGND VPWR VPWR U$$81/X sky130_fd_sc_hd__xor2_1
XU$$92 U$$92/A1 U$$96/A2 U$$94/A1 U$$96/B2 VGND VGND VPWR VPWR U$$93/A sky130_fd_sc_hd__a22o_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_107_1 U$$3812/X U$$3945/X U$$4078/X VGND VGND VPWR VPWR dadda_fa_4_108_0/CIN
+ dadda_fa_4_107_2/A sky130_fd_sc_hd__fa_1
XFILLER_106_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_48_3 dadda_fa_3_48_3/A dadda_fa_3_48_3/B dadda_fa_3_48_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_1/B dadda_fa_4_48_2/CIN sky130_fd_sc_hd__fa_1
XU$$1204 U$$930/A1 U$$1230/A2 U$$932/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1205/A sky130_fd_sc_hd__a22o_1
XFILLER_55_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1215 U$$1215/A U$$1221/B VGND VGND VPWR VPWR U$$1215/X sky130_fd_sc_hd__xor2_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1226 U$$678/A1 U$$1226/A2 U$$678/B1 U$$1226/B2 VGND VGND VPWR VPWR U$$1227/A sky130_fd_sc_hd__a22o_1
XU$$1237 U$$1235/Y input10/X U$$1233/A U$$1236/X U$$1233/Y VGND VGND VPWR VPWR U$$1237/X
+ sky130_fd_sc_hd__a32o_2
XU$$1248 U$$1248/A U$$1282/B VGND VGND VPWR VPWR U$$1248/X sky130_fd_sc_hd__xor2_1
XFILLER_44_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1259 U$$983/B1 U$$1295/A2 U$$850/A1 U$$1295/B2 VGND VGND VPWR VPWR U$$1260/A sky130_fd_sc_hd__a22o_1
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1031 final_adder.U$$7/SUM final_adder.U$$1031/B VGND VGND VPWR VPWR
+ output362/A sky130_fd_sc_hd__xor2_1
XFILLER_144_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1042 final_adder.U$$236/A final_adder.U$$737/X VGND VGND VPWR VPWR
+ output294/A sky130_fd_sc_hd__xor2_1
XFILLER_7_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1053 final_adder.U$$226/B final_adder.U$$997/X VGND VGND VPWR VPWR
+ output306/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1064 final_adder.U$$214/A final_adder.U$$827/X VGND VGND VPWR VPWR
+ output319/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1075 final_adder.U$$204/B final_adder.U$$975/X VGND VGND VPWR VPWR
+ output331/A sky130_fd_sc_hd__xor2_1
XU$$4439_1867 VGND VGND VPWR VPWR U$$4439_1867/HI U$$4439/B sky130_fd_sc_hd__conb_1
XFILLER_172_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1086 final_adder.U$$192/A final_adder.U$$805/X VGND VGND VPWR VPWR
+ output343/A sky130_fd_sc_hd__xor2_1
XFILLER_109_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1097 final_adder.U$$182/B final_adder.U$$953/X VGND VGND VPWR VPWR
+ output355/A sky130_fd_sc_hd__xor2_1
XFILLER_139_1040 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1360 fanout1364/X VGND VGND VPWR VPWR U$$3258/B sky130_fd_sc_hd__clkbuf_4
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_50_3 dadda_fa_2_50_3/A dadda_fa_2_50_3/B dadda_fa_2_50_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_1/B dadda_fa_3_50_3/B sky130_fd_sc_hd__fa_1
Xfanout1371 U$$3119/B VGND VGND VPWR VPWR U$$3147/B sky130_fd_sc_hd__clkbuf_4
XFILLER_66_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1382 input38/X VGND VGND VPWR VPWR U$$2990/B sky130_fd_sc_hd__buf_6
Xfanout1393 U$$260/B VGND VGND VPWR VPWR U$$220/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_43_2 U$$2753/X U$$2886/X input194/X VGND VGND VPWR VPWR dadda_fa_3_44_1/A
+ dadda_fa_3_43_3/A sky130_fd_sc_hd__fa_1
XU$$3140 U$$3960/B1 U$$3148/A2 U$$3825/B1 U$$3148/B2 VGND VGND VPWR VPWR U$$3141/A
+ sky130_fd_sc_hd__a22o_1
XU$$3151 U$$3151/A VGND VGND VPWR VPWR U$$3151/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_5_20_1 dadda_fa_5_20_1/A dadda_fa_5_20_1/B dadda_fa_5_20_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_21_0/B dadda_fa_7_20_0/A sky130_fd_sc_hd__fa_1
XU$$3162 U$$3162/A U$$3196/B VGND VGND VPWR VPWR U$$3162/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_36_1 U$$1143/X U$$1276/X U$$1409/X VGND VGND VPWR VPWR dadda_fa_3_37_0/CIN
+ dadda_fa_3_36_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3173 U$$4406/A1 U$$3257/A2 U$$4408/A1 U$$3257/B2 VGND VGND VPWR VPWR U$$3174/A
+ sky130_fd_sc_hd__a22o_1
XU$$3184 U$$3184/A U$$3208/B VGND VGND VPWR VPWR U$$3184/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_13_0 dadda_fa_5_13_0/A dadda_fa_5_13_0/B dadda_fa_5_13_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_14_0/A dadda_fa_6_13_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_34_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3195 U$$4428/A1 U$$3199/A2 U$$4430/A1 U$$3199/B2 VGND VGND VPWR VPWR U$$3196/A
+ sky130_fd_sc_hd__a22o_1
XU$$2450 U$$2450/A U$$2456/B VGND VGND VPWR VPWR U$$2450/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_29_0 U$$65/X U$$198/X U$$331/X VGND VGND VPWR VPWR dadda_fa_3_30_1/B dadda_fa_3_29_3/A
+ sky130_fd_sc_hd__fa_1
XFILLER_50_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2461 U$$954/A1 U$$2463/A2 U$$956/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2462/A sky130_fd_sc_hd__a22o_1
XU$$2472 U$$2472/A1 U$$2548/A2 U$$828/B1 U$$2548/B2 VGND VGND VPWR VPWR U$$2473/A
+ sky130_fd_sc_hd__a22o_1
XU$$2483 U$$2483/A U$$2541/B VGND VGND VPWR VPWR U$$2483/X sky130_fd_sc_hd__xor2_1
XU$$2494 U$$2631/A1 U$$2532/A2 U$$2631/B1 U$$2532/B2 VGND VGND VPWR VPWR U$$2495/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1760 U$$2443/B1 U$$1760/A2 U$$2310/A1 U$$1760/B2 VGND VGND VPWR VPWR U$$1761/A
+ sky130_fd_sc_hd__a22o_1
XU$$1771 U$$1771/A U$$1777/B VGND VGND VPWR VPWR U$$1771/X sky130_fd_sc_hd__xor2_1
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1782 input19/X VGND VGND VPWR VPWR U$$1784/B sky130_fd_sc_hd__inv_1
XU$$1793 U$$2887/B1 U$$1829/A2 U$$2754/A1 U$$1829/B2 VGND VGND VPWR VPWR U$$1794/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput70 b[14] VGND VGND VPWR VPWR input70/X sky130_fd_sc_hd__clkbuf_4
Xinput81 b[24] VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__buf_4
XFILLER_116_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput92 b[34] VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_58_2 dadda_fa_4_58_2/A dadda_fa_4_58_2/B dadda_fa_4_58_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_59_0/CIN dadda_fa_5_58_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$401 final_adder.U$$400/B final_adder.U$$279/X final_adder.U$$275/X
+ VGND VGND VPWR VPWR final_adder.U$$401/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$412 final_adder.U$$416/B final_adder.U$$412/B VGND VGND VPWR VPWR
+ final_adder.U$$536/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$423 final_adder.U$$422/B final_adder.U$$301/X final_adder.U$$297/X
+ VGND VGND VPWR VPWR final_adder.U$$423/X sky130_fd_sc_hd__a21o_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$434 final_adder.U$$438/B final_adder.U$$434/B VGND VGND VPWR VPWR
+ final_adder.U$$558/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$445 final_adder.U$$444/B final_adder.U$$323/X final_adder.U$$319/X
+ VGND VGND VPWR VPWR final_adder.U$$445/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$456 final_adder.U$$460/B final_adder.U$$456/B VGND VGND VPWR VPWR
+ final_adder.U$$580/B sky130_fd_sc_hd__and2_1
Xdadda_fa_7_28_0 dadda_fa_7_28_0/A dadda_fa_7_28_0/B dadda_fa_7_28_0/CIN VGND VGND
+ VPWR VPWR _325_/D _196_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$467 final_adder.U$$466/B final_adder.U$$345/X final_adder.U$$341/X
+ VGND VGND VPWR VPWR final_adder.U$$467/X sky130_fd_sc_hd__a21o_1
XU$$306 U$$443/A1 U$$338/A2 U$$34/A1 U$$338/B2 VGND VGND VPWR VPWR U$$307/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$478 final_adder.U$$482/B final_adder.U$$478/B VGND VGND VPWR VPWR
+ final_adder.U$$602/B sky130_fd_sc_hd__and2_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$317 U$$317/A U$$339/B VGND VGND VPWR VPWR U$$317/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$489 final_adder.U$$488/B final_adder.U$$367/X final_adder.U$$363/X
+ VGND VGND VPWR VPWR final_adder.U$$489/X sky130_fd_sc_hd__a21o_1
XFILLER_26_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$328 U$$465/A1 U$$362/A2 U$$465/B1 U$$362/B2 VGND VGND VPWR VPWR U$$329/A sky130_fd_sc_hd__a22o_1
XU$$339 U$$339/A U$$339/B VGND VGND VPWR VPWR U$$339/X sky130_fd_sc_hd__xor2_1
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1000 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_102_0_1932 VGND VGND VPWR VPWR dadda_fa_2_102_0/A dadda_fa_2_102_0_1932/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_60_2 dadda_fa_3_60_2/A dadda_fa_3_60_2/B dadda_fa_3_60_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_1/A dadda_fa_4_60_2/B sky130_fd_sc_hd__fa_1
XFILLER_0_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_53_1 dadda_fa_3_53_1/A dadda_fa_3_53_1/B dadda_fa_3_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_0/CIN dadda_fa_4_53_2/A sky130_fd_sc_hd__fa_1
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_69_1 U$$810/X U$$943/X U$$1076/X VGND VGND VPWR VPWR dadda_fa_1_70_6/B
+ dadda_fa_1_69_8/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_30_0 dadda_fa_6_30_0/A dadda_fa_6_30_0/B dadda_fa_6_30_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_31_0/B dadda_fa_7_30_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_46_0 dadda_fa_3_46_0/A dadda_fa_3_46_0/B dadda_fa_3_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_0/B dadda_fa_4_46_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_91_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$840 U$$840/A1 U$$876/A2 U$$840/B1 U$$876/B2 VGND VGND VPWR VPWR U$$841/A sky130_fd_sc_hd__a22o_1
XU$$851 U$$851/A U$$895/B VGND VGND VPWR VPWR U$$851/X sky130_fd_sc_hd__xor2_1
XU$$862 U$$997/B1 U$$898/A2 U$$864/A1 U$$898/B2 VGND VGND VPWR VPWR U$$863/A sky130_fd_sc_hd__a22o_1
XU$$1001 U$$999/B1 U$$981/A2 U$$866/A1 U$$981/B2 VGND VGND VPWR VPWR U$$1002/A sky130_fd_sc_hd__a22o_1
XU$$1012 U$$1012/A U$$1046/B VGND VGND VPWR VPWR U$$1012/X sky130_fd_sc_hd__xor2_1
XU$$873 U$$873/A U$$875/B VGND VGND VPWR VPWR U$$873/X sky130_fd_sc_hd__xor2_1
XU$$1023 U$$64/A1 U$$997/A2 U$$64/B1 U$$997/B2 VGND VGND VPWR VPWR U$$1024/A sky130_fd_sc_hd__a22o_1
XU$$884 U$$884/A1 U$$902/A2 U$$884/B1 U$$902/B2 VGND VGND VPWR VPWR U$$885/A sky130_fd_sc_hd__a22o_1
XFILLER_90_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$895 U$$895/A U$$895/B VGND VGND VPWR VPWR U$$895/X sky130_fd_sc_hd__xor2_1
XU$$1034 U$$1034/A U$$1062/B VGND VGND VPWR VPWR U$$1034/X sky130_fd_sc_hd__xor2_1
XFILLER_31_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1045 U$$906/B1 U$$1087/A2 U$$773/A1 U$$1087/B2 VGND VGND VPWR VPWR U$$1046/A sky130_fd_sc_hd__a22o_1
XU$$1056 U$$1056/A U$$990/B VGND VGND VPWR VPWR U$$1056/X sky130_fd_sc_hd__xor2_1
XU$$1067 U$$930/A1 U$$1075/A2 U$$932/A1 U$$1075/B2 VGND VGND VPWR VPWR U$$1068/A sky130_fd_sc_hd__a22o_1
XU$$1078 U$$1078/A U$$1094/B VGND VGND VPWR VPWR U$$1078/X sky130_fd_sc_hd__xor2_1
XU$$1089 U$$952/A1 U$$1093/A2 U$$954/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1090/A sky130_fd_sc_hd__a22o_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_103_0 dadda_fa_7_103_0/A dadda_fa_7_103_0/B dadda_fa_7_103_0/CIN VGND
+ VGND VPWR VPWR _400_/D _271_/D sky130_fd_sc_hd__fa_1
XFILLER_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_98_3 U$$3528/X U$$3661/X U$$3794/X VGND VGND VPWR VPWR dadda_fa_3_99_1/CIN
+ dadda_fa_3_98_3/B sky130_fd_sc_hd__fa_1
XFILLER_160_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_5_68_1 dadda_fa_5_68_1/A dadda_fa_5_68_1/B dadda_fa_5_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_69_0/B dadda_fa_7_68_0/A sky130_fd_sc_hd__fa_1
Xfanout608 U$$1758/A2 VGND VGND VPWR VPWR U$$1774/A2 sky130_fd_sc_hd__buf_4
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout619 U$$1621/A2 VGND VGND VPWR VPWR U$$1625/A2 sky130_fd_sc_hd__buf_6
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1190 U$$3048/B1 VGND VGND VPWR VPWR U$$447/A1 sky130_fd_sc_hd__buf_4
XFILLER_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_107_0 U$$3013/Y U$$3147/X U$$3280/X VGND VGND VPWR VPWR dadda_fa_3_108_3/CIN
+ dadda_fa_4_107_0/A sky130_fd_sc_hd__fa_1
XU$$2280 U$$773/A1 U$$2282/A2 U$$773/B1 U$$2282/B2 VGND VGND VPWR VPWR U$$2281/A sky130_fd_sc_hd__a22o_1
XU$$2291 U$$2291/A U$$2327/B VGND VGND VPWR VPWR U$$2291/X sky130_fd_sc_hd__xor2_1
XFILLER_167_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1590 U$$1590/A U$$1594/B VGND VGND VPWR VPWR U$$1590/X sky130_fd_sc_hd__xor2_1
XFILLER_139_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_70_1 dadda_fa_4_70_1/A dadda_fa_4_70_1/B dadda_fa_4_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_71_0/B dadda_fa_5_70_1/B sky130_fd_sc_hd__fa_1
XFILLER_116_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_86_1 U$$1908/X U$$2041/X U$$2174/X VGND VGND VPWR VPWR dadda_fa_2_87_3/A
+ dadda_fa_2_86_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_63_0 dadda_fa_4_63_0/A dadda_fa_4_63_0/B dadda_fa_4_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_64_0/A dadda_fa_5_63_1/A sky130_fd_sc_hd__fa_1
XFILLER_77_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_79_0 U$$1095/Y U$$1229/X U$$1362/X VGND VGND VPWR VPWR dadda_fa_2_80_0/B
+ dadda_fa_2_79_3/B sky130_fd_sc_hd__fa_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$220 final_adder.U$$220/A final_adder.U$$220/B VGND VGND VPWR VPWR
+ final_adder.U$$348/B sky130_fd_sc_hd__and2_1
XFILLER_40_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$231 final_adder.U$$230/B final_adder.U$$231/A2 final_adder.U$$231/B1
+ VGND VGND VPWR VPWR final_adder.U$$231/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$242 final_adder.U$$242/A final_adder.U$$242/B VGND VGND VPWR VPWR
+ final_adder.U$$370/B sky130_fd_sc_hd__and2_1
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3909 U$$3909/A U$$3973/A VGND VGND VPWR VPWR U$$3909/X sky130_fd_sc_hd__xor2_1
XFILLER_94_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$253 final_adder.U$$3/SUM final_adder.U$$253/A2 final_adder.U$$3/COUT
+ VGND VGND VPWR VPWR final_adder.U$$253/X sky130_fd_sc_hd__a21o_1
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$264 final_adder.U$$266/B final_adder.U$$264/B VGND VGND VPWR VPWR
+ final_adder.U$$390/B sky130_fd_sc_hd__and2_1
XFILLER_27_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$103 U$$103/A U$$99/B VGND VGND VPWR VPWR U$$103/X sky130_fd_sc_hd__xor2_1
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$275 final_adder.U$$274/B final_adder.U$$149/X final_adder.U$$147/X
+ VGND VGND VPWR VPWR final_adder.U$$275/X sky130_fd_sc_hd__a21o_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$114 U$$386/B1 U$$120/A2 U$$253/A1 U$$120/B2 VGND VGND VPWR VPWR U$$115/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$286 final_adder.U$$288/B final_adder.U$$286/B VGND VGND VPWR VPWR
+ final_adder.U$$412/B sky130_fd_sc_hd__and2_1
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$125 U$$125/A U$$3/A VGND VGND VPWR VPWR U$$125/X sky130_fd_sc_hd__xor2_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$297 final_adder.U$$296/B final_adder.U$$171/X final_adder.U$$169/X
+ VGND VGND VPWR VPWR final_adder.U$$297/X sky130_fd_sc_hd__a21o_1
XU$$136 U$$99/B VGND VGND VPWR VPWR U$$136/Y sky130_fd_sc_hd__inv_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$147 U$$10/A1 U$$179/A2 U$$12/A1 U$$179/B2 VGND VGND VPWR VPWR U$$148/A sky130_fd_sc_hd__a22o_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$158 U$$158/A U$$180/B VGND VGND VPWR VPWR U$$158/X sky130_fd_sc_hd__xor2_1
XU$$169 U$$443/A1 U$$207/A2 U$$34/A1 U$$207/B2 VGND VGND VPWR VPWR U$$170/A sky130_fd_sc_hd__a22o_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_393_ _397_/CLK _393_/D VGND VGND VPWR VPWR _393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_78_0 dadda_fa_6_78_0/A dadda_fa_6_78_0/B dadda_fa_6_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_79_0/B dadda_fa_7_78_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$670 U$$805/B1 U$$674/A2 U$$672/A1 U$$674/B2 VGND VGND VPWR VPWR U$$671/A sky130_fd_sc_hd__a22o_1
XFILLER_91_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$681 U$$681/A U$$684/A VGND VGND VPWR VPWR U$$681/X sky130_fd_sc_hd__xor2_1
XU$$692 U$$692/A U$$744/B VGND VGND VPWR VPWR U$$692/X sky130_fd_sc_hd__xor2_1
XFILLER_17_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_80_0 dadda_fa_5_80_0/A dadda_fa_5_80_0/B dadda_fa_5_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_81_0/A dadda_fa_6_80_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_96_0 U$$2460/X U$$2593/X U$$2726/X VGND VGND VPWR VPWR dadda_fa_3_97_0/B
+ dadda_fa_3_96_2/B sky130_fd_sc_hd__fa_1
XFILLER_144_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout405 U$$819/A2 VGND VGND VPWR VPWR U$$771/A2 sky130_fd_sc_hd__buf_4
Xfanout416 U$$4289/A2 VGND VGND VPWR VPWR U$$4295/A2 sky130_fd_sc_hd__buf_4
Xfanout427 U$$543/A2 VGND VGND VPWR VPWR U$$539/A2 sky130_fd_sc_hd__buf_4
XFILLER_59_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_72_7 dadda_fa_1_72_7/A dadda_fa_1_72_7/B dadda_fa_1_72_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_73_2/CIN dadda_fa_2_72_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_98_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout438 U$$4190/A2 VGND VGND VPWR VPWR U$$4224/A2 sky130_fd_sc_hd__buf_4
Xfanout449 U$$4/X VGND VGND VPWR VPWR U$$102/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_65_6 dadda_fa_1_65_6/A dadda_fa_1_65_6/B dadda_fa_1_65_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_66_2/B dadda_fa_2_65_5/B sky130_fd_sc_hd__fa_1
XFILLER_104_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_58_5 U$$3581/X U$$3714/X U$$3847/X VGND VGND VPWR VPWR dadda_fa_2_59_2/A
+ dadda_fa_2_58_5/A sky130_fd_sc_hd__fa_1
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_95_0 dadda_fa_7_95_0/A dadda_fa_7_95_0/B dadda_fa_7_95_0/CIN VGND VGND
+ VPWR VPWR _392_/D _263_/D sky130_fd_sc_hd__fa_1
XFILLER_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout950 fanout957/X VGND VGND VPWR VPWR U$$86/A1 sky130_fd_sc_hd__buf_4
Xfanout961 fanout966/X VGND VGND VPWR VPWR U$$3509/A1 sky130_fd_sc_hd__buf_6
XU$$4407 U$$4407/A U$$4407/B VGND VGND VPWR VPWR U$$4407/X sky130_fd_sc_hd__xor2_1
Xfanout972 fanout975/X VGND VGND VPWR VPWR U$$80/B1 sky130_fd_sc_hd__buf_2
XU$$4418 input69/X U$$4388/X input70/X U$$4508/B2 VGND VGND VPWR VPWR U$$4419/A sky130_fd_sc_hd__a22o_1
XU$$4429 U$$4429/A U$$4429/B VGND VGND VPWR VPWR U$$4429/X sky130_fd_sc_hd__xor2_1
Xfanout983 fanout984/X VGND VGND VPWR VPWR U$$4464/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout994 fanout999/A VGND VGND VPWR VPWR U$$898/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_6_110_0 dadda_fa_6_110_0/A dadda_fa_6_110_0/B dadda_fa_6_110_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_111_0/B dadda_fa_7_110_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3706 U$$3706/A U$$3790/B VGND VGND VPWR VPWR U$$3706/X sky130_fd_sc_hd__xor2_1
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3717 U$$4400/B1 U$$3757/A2 U$$4265/B1 U$$3757/B2 VGND VGND VPWR VPWR U$$3718/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3728 U$$3728/A U$$3734/B VGND VGND VPWR VPWR U$$3728/X sky130_fd_sc_hd__xor2_1
XFILLER_45_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3739 U$$4150/A1 U$$3739/A2 U$$4152/A1 U$$3739/B2 VGND VGND VPWR VPWR U$$3740/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_3 dadda_fa_3_30_3/A dadda_fa_3_30_3/B dadda_fa_3_30_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_31_1/B dadda_fa_4_30_2/CIN sky130_fd_sc_hd__fa_1
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_23_2 U$$1117/X U$$1250/X U$$1383/X VGND VGND VPWR VPWR dadda_fa_4_24_1/A
+ dadda_fa_4_23_2/B sky130_fd_sc_hd__fa_1
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_376_ _397_/CLK _376_/D VGND VGND VPWR VPWR _376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1093_1781 VGND VGND VPWR VPWR U$$1093_1781/HI U$$1093/B1 sky130_fd_sc_hd__conb_1
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_75_5 dadda_fa_2_75_5/A dadda_fa_2_75_5/B dadda_fa_2_75_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_2/A dadda_fa_4_75_0/A sky130_fd_sc_hd__fa_1
XFILLER_68_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_68_4 dadda_fa_2_68_4/A dadda_fa_2_68_4/B dadda_fa_2_68_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_1/CIN dadda_fa_3_68_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_105_1 dadda_fa_5_105_1/A dadda_fa_5_105_1/B dadda_fa_5_105_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_106_0/B dadda_fa_7_105_0/A sky130_fd_sc_hd__fa_1
XFILLER_105_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_70_4 U$$3871/X U$$4004/X U$$4137/X VGND VGND VPWR VPWR dadda_fa_2_71_1/CIN
+ dadda_fa_2_70_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_101_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_63_3 U$$3591/X U$$3724/X U$$3857/X VGND VGND VPWR VPWR dadda_fa_2_64_1/B
+ dadda_fa_2_63_4/B sky130_fd_sc_hd__fa_1
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_40_2 dadda_fa_4_40_2/A dadda_fa_4_40_2/B dadda_fa_4_40_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_41_0/CIN dadda_fa_5_40_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_56_2 U$$1981/X U$$2114/X U$$2247/X VGND VGND VPWR VPWR dadda_fa_2_57_1/A
+ dadda_fa_2_56_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_33_1 dadda_fa_4_33_1/A dadda_fa_4_33_1/B dadda_fa_4_33_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_34_0/B dadda_fa_5_33_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_49_1 U$$504/X U$$637/X U$$770/X VGND VGND VPWR VPWR dadda_fa_2_50_1/A
+ dadda_fa_2_49_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_7_10_0 dadda_fa_7_10_0/A dadda_fa_7_10_0/B dadda_fa_7_10_0/CIN VGND VGND
+ VPWR VPWR _307_/D _178_/D sky130_fd_sc_hd__fa_1
XFILLER_43_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_26_0 dadda_fa_4_26_0/A dadda_fa_4_26_0/B dadda_fa_4_26_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_27_0/A dadda_fa_5_26_1/A sky130_fd_sc_hd__fa_1
XFILLER_70_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_230_ _359_/CLK _230_/D VGND VGND VPWR VPWR _230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_78_3 dadda_fa_3_78_3/A dadda_fa_3_78_3/B dadda_fa_3_78_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_1/B dadda_fa_4_78_2/CIN sky130_fd_sc_hd__fa_1
Xfanout1701 U$$2844/B1 VGND VGND VPWR VPWR U$$2707/B1 sky130_fd_sc_hd__buf_4
Xfanout1712 fanout1718/X VGND VGND VPWR VPWR U$$2979/B1 sky130_fd_sc_hd__buf_4
XFILLER_151_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1723 input106/X VGND VGND VPWR VPWR U$$650/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_172_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1734 input105/X VGND VGND VPWR VPWR U$$3249/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout1745 U$$505/B1 VGND VGND VPWR VPWR U$$2973/A1 sky130_fd_sc_hd__buf_4
Xfanout1756 input102/X VGND VGND VPWR VPWR U$$3243/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_77_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4204 U$$4341/A1 U$$4226/A2 U$$4480/A1 U$$4226/B2 VGND VGND VPWR VPWR U$$4205/A
+ sky130_fd_sc_hd__a22o_1
XU$$4215 U$$4215/A U$$4215/B VGND VGND VPWR VPWR U$$4215/X sky130_fd_sc_hd__xor2_1
Xfanout1767 U$$3515/B1 VGND VGND VPWR VPWR U$$4476/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout780 U$$2977/B2 VGND VGND VPWR VPWR U$$2937/B2 sky130_fd_sc_hd__buf_6
XU$$4226 U$$4226/A1 U$$4226/A2 U$$4226/B1 U$$4226/B2 VGND VGND VPWR VPWR U$$4227/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1778 U$$912/A1 VGND VGND VPWR VPWR U$$3650/B1 sky130_fd_sc_hd__buf_6
Xfanout791 U$$340/B2 VGND VGND VPWR VPWR U$$312/B2 sky130_fd_sc_hd__buf_2
XU$$4237 U$$4237/A U$$4241/B VGND VGND VPWR VPWR U$$4237/X sky130_fd_sc_hd__xor2_1
XU$$3503 U$$3638/B1 U$$3505/A2 U$$3503/B1 U$$3505/B2 VGND VGND VPWR VPWR U$$3504/A
+ sky130_fd_sc_hd__a22o_1
XU$$4248 input59/X VGND VGND VPWR VPWR U$$4250/B sky130_fd_sc_hd__inv_1
Xdadda_ha_3_15_0 U$$37/X U$$170/X VGND VGND VPWR VPWR dadda_fa_4_16_2/A dadda_ha_3_15_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$4259 U$$4396/A1 U$$4295/A2 U$$4259/B1 U$$4295/B2 VGND VGND VPWR VPWR U$$4260/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3514 U$$3514/A U$$3558/B VGND VGND VPWR VPWR U$$3514/X sky130_fd_sc_hd__xor2_1
XU$$3525 U$$4482/B1 U$$3549/A2 U$$4349/A1 U$$3549/B2 VGND VGND VPWR VPWR U$$3526/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3536 U$$3536/A U$$3548/B VGND VGND VPWR VPWR U$$3536/X sky130_fd_sc_hd__xor2_1
XU$$2802 U$$4309/A1 U$$2844/A2 U$$3763/A1 U$$2844/B2 VGND VGND VPWR VPWR U$$2803/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3547 U$$3684/A1 U$$3549/A2 U$$3684/B1 U$$3549/B2 VGND VGND VPWR VPWR U$$3548/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3558 U$$3558/A U$$3558/B VGND VGND VPWR VPWR U$$3558/X sky130_fd_sc_hd__xor2_1
XU$$2813 U$$2813/A U$$2873/B VGND VGND VPWR VPWR U$$2813/X sky130_fd_sc_hd__xor2_1
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2824 U$$3509/A1 U$$2840/A2 U$$3509/B1 U$$2840/B2 VGND VGND VPWR VPWR U$$2825/A
+ sky130_fd_sc_hd__a22o_1
XU$$3569 U$$3569/A U$$3615/B VGND VGND VPWR VPWR U$$3569/X sky130_fd_sc_hd__xor2_1
XU$$2835 U$$2835/A U$$2841/B VGND VGND VPWR VPWR U$$2835/X sky130_fd_sc_hd__xor2_1
XFILLER_65_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2846 U$$4353/A1 U$$2874/A2 U$$4353/B1 U$$2874/B2 VGND VGND VPWR VPWR U$$2847/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2857 U$$2857/A U$$2873/B VGND VGND VPWR VPWR U$$2857/X sky130_fd_sc_hd__xor2_1
XFILLER_34_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2868 U$$3416/A1 U$$2872/A2 U$$3418/A1 U$$2872/B2 VGND VGND VPWR VPWR U$$2869/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2879 U$$2974/B VGND VGND VPWR VPWR U$$2879/Y sky130_fd_sc_hd__inv_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_359_ _359_/CLK _359_/D VGND VGND VPWR VPWR _359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_80_3 dadda_fa_2_80_3/A dadda_fa_2_80_3/B dadda_fa_2_80_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_1/B dadda_fa_3_80_3/B sky130_fd_sc_hd__fa_1
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_73_2 dadda_fa_2_73_2/A dadda_fa_2_73_2/B dadda_fa_2_73_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_1/A dadda_fa_3_73_3/A sky130_fd_sc_hd__fa_1
XFILLER_130_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_50_1 dadda_fa_5_50_1/A dadda_fa_5_50_1/B dadda_fa_5_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_51_0/B dadda_fa_7_50_0/A sky130_fd_sc_hd__fa_1
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_66_1 dadda_fa_2_66_1/A dadda_fa_2_66_1/B dadda_fa_2_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_0/CIN dadda_fa_3_66_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$819 final_adder.U$$786/A final_adder.U$$619/X final_adder.U$$707/X
+ VGND VGND VPWR VPWR final_adder.U$$819/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_5_43_0 dadda_fa_5_43_0/A dadda_fa_5_43_0/B dadda_fa_5_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_44_0/A dadda_fa_6_43_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_59_0 dadda_fa_2_59_0/A dadda_fa_2_59_0/B dadda_fa_2_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_0/B dadda_fa_3_59_2/B sky130_fd_sc_hd__fa_1
XFILLER_111_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput2 a[10] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$0 _296_/Q _168_/Q VGND VGND VPWR VPWR final_adder.U$$255/A2 final_adder.U$$0/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_69_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_88_2 dadda_fa_4_88_2/A dadda_fa_4_88_2/B dadda_fa_4_88_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_89_0/CIN dadda_fa_5_88_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4391_1843 VGND VGND VPWR VPWR U$$4391_1843/HI U$$4391/B sky130_fd_sc_hd__conb_1
Xoutput350 output350/A VGND VGND VPWR VPWR o[69] sky130_fd_sc_hd__buf_2
Xoutput361 output361/A VGND VGND VPWR VPWR o[79] sky130_fd_sc_hd__buf_2
XFILLER_160_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_58_0 dadda_fa_7_58_0/A dadda_fa_7_58_0/B dadda_fa_7_58_0/CIN VGND VGND
+ VPWR VPWR _355_/D _226_/D sky130_fd_sc_hd__fa_1
Xoutput372 output372/A VGND VGND VPWR VPWR o[89] sky130_fd_sc_hd__buf_2
XFILLER_0_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput383 output383/A VGND VGND VPWR VPWR o[99] sky130_fd_sc_hd__buf_2
XFILLER_86_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1008 fanout1011/X VGND VGND VPWR VPWR U$$3908/B1 sky130_fd_sc_hd__buf_2
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1019 input90/X VGND VGND VPWR VPWR U$$4182/A1 sky130_fd_sc_hd__buf_6
XFILLER_126_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_0 U$$1991/X U$$2124/X U$$2257/X VGND VGND VPWR VPWR dadda_fa_2_62_0/B
+ dadda_fa_2_61_3/B sky130_fd_sc_hd__fa_1
XFILLER_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2109 U$$876/A1 U$$2147/A2 U$$878/A1 U$$2147/B2 VGND VGND VPWR VPWR U$$2110/A sky130_fd_sc_hd__a22o_1
XFILLER_83_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1408 U$$447/B1 U$$1414/A2 U$$314/A1 U$$1414/B2 VGND VGND VPWR VPWR U$$1409/A sky130_fd_sc_hd__a22o_1
XU$$1419 U$$1419/A U$$1433/B VGND VGND VPWR VPWR U$$1419/X sky130_fd_sc_hd__xor2_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_213_ _342_/CLK _213_/D VGND VGND VPWR VPWR _213_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_169_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_90_2 dadda_fa_3_90_2/A dadda_fa_3_90_2/B dadda_fa_3_90_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_1/A dadda_fa_4_90_2/B sky130_fd_sc_hd__fa_1
XFILLER_136_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_83_1 dadda_fa_3_83_1/A dadda_fa_3_83_1/B dadda_fa_3_83_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_0/CIN dadda_fa_4_83_2/A sky130_fd_sc_hd__fa_1
XFILLER_83_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_60_0 dadda_fa_6_60_0/A dadda_fa_6_60_0/B dadda_fa_6_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_61_0/B dadda_fa_7_60_0/CIN sky130_fd_sc_hd__fa_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_76_0 dadda_fa_3_76_0/A dadda_fa_3_76_0/B dadda_fa_3_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_0/B dadda_fa_4_76_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1520 U$$3447/B1 VGND VGND VPWR VPWR U$$24/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1531 U$$2897/A1 VGND VGND VPWR VPWR U$$2758/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1542 input124/X VGND VGND VPWR VPWR U$$956/A1 sky130_fd_sc_hd__buf_4
Xfanout1553 U$$3692/B1 VGND VGND VPWR VPWR U$$3418/B1 sky130_fd_sc_hd__buf_4
XU$$4001 U$$987/A1 U$$4005/A2 U$$4001/B1 U$$4005/B2 VGND VGND VPWR VPWR U$$4002/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1564 input122/X VGND VGND VPWR VPWR U$$4514/A1 sky130_fd_sc_hd__buf_4
XU$$4012 U$$4012/A U$$4058/B VGND VGND VPWR VPWR U$$4012/X sky130_fd_sc_hd__xor2_1
XU$$4023 U$$4295/B1 U$$4045/A2 U$$4436/A1 U$$4045/B2 VGND VGND VPWR VPWR U$$4024/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1575 U$$4402/A1 VGND VGND VPWR VPWR U$$3030/B1 sky130_fd_sc_hd__buf_4
XFILLER_66_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4034 U$$4034/A U$$4040/B VGND VGND VPWR VPWR U$$4034/X sky130_fd_sc_hd__xor2_1
Xfanout1586 input12/X VGND VGND VPWR VPWR U$$127/B sky130_fd_sc_hd__buf_6
XFILLER_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3300 U$$4257/B1 U$$3340/A2 U$$4259/B1 U$$3340/B2 VGND VGND VPWR VPWR U$$3301/A
+ sky130_fd_sc_hd__a22o_1
XU$$4045 U$$4456/A1 U$$4045/A2 U$$4458/A1 U$$4045/B2 VGND VGND VPWR VPWR U$$4046/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1597 U$$2729/A1 VGND VGND VPWR VPWR U$$4234/B1 sky130_fd_sc_hd__clkbuf_4
XU$$3311 U$$3311/A U$$3349/B VGND VGND VPWR VPWR U$$3311/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_112_1 dadda_fa_4_112_1/A dadda_fa_4_112_1/B dadda_fa_4_112_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_113_0/B dadda_fa_5_112_1/B sky130_fd_sc_hd__fa_1
XU$$4056 U$$4056/A U$$4058/B VGND VGND VPWR VPWR U$$4056/X sky130_fd_sc_hd__xor2_1
XU$$3322 U$$3870/A1 U$$3338/A2 U$$3322/B1 U$$3338/B2 VGND VGND VPWR VPWR U$$3323/A
+ sky130_fd_sc_hd__a22o_1
XU$$4067 U$$4341/A1 U$$4093/A2 U$$4480/A1 U$$4093/B2 VGND VGND VPWR VPWR U$$4068/A
+ sky130_fd_sc_hd__a22o_1
XU$$3333 U$$3333/A U$$3373/B VGND VGND VPWR VPWR U$$3333/X sky130_fd_sc_hd__xor2_1
XU$$4078 U$$4078/A U$$4082/B VGND VGND VPWR VPWR U$$4078/X sky130_fd_sc_hd__xor2_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4089 U$$4226/A1 U$$4107/A2 U$$4226/B1 U$$4107/B2 VGND VGND VPWR VPWR U$$4090/A
+ sky130_fd_sc_hd__a22o_1
XU$$3344 U$$878/A1 U$$3390/A2 U$$878/B1 U$$3390/B2 VGND VGND VPWR VPWR U$$3345/A sky130_fd_sc_hd__a22o_1
XU$$3355 U$$3355/A U$$3425/A VGND VGND VPWR VPWR U$$3355/X sky130_fd_sc_hd__xor2_1
XU$$2610 U$$2610/A U$$2678/B VGND VGND VPWR VPWR U$$2610/X sky130_fd_sc_hd__xor2_1
XU$$2621 U$$2758/A1 U$$2665/A2 U$$2758/B1 U$$2665/B2 VGND VGND VPWR VPWR U$$2622/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_38_5 dadda_fa_2_38_5/A dadda_fa_2_38_5/B dadda_fa_2_38_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_39_2/A dadda_fa_4_38_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_4_105_0 dadda_fa_4_105_0/A dadda_fa_4_105_0/B dadda_fa_4_105_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_106_0/A dadda_fa_5_105_1/A sky130_fd_sc_hd__fa_1
XU$$3366 U$$3638/B1 U$$3372/A2 U$$3503/B1 U$$3372/B2 VGND VGND VPWR VPWR U$$3367/A
+ sky130_fd_sc_hd__a22o_1
XU$$3377 U$$3377/A U$$3425/A VGND VGND VPWR VPWR U$$3377/X sky130_fd_sc_hd__xor2_1
XU$$2632 U$$2632/A U$$2668/B VGND VGND VPWR VPWR U$$2632/X sky130_fd_sc_hd__xor2_1
XFILLER_80_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2643 U$$4150/A1 U$$2681/A2 U$$4152/A1 U$$2681/B2 VGND VGND VPWR VPWR U$$2644/A
+ sky130_fd_sc_hd__a22o_1
XU$$3388 U$$920/B1 U$$3390/A2 U$$787/A1 U$$3390/B2 VGND VGND VPWR VPWR U$$3389/A sky130_fd_sc_hd__a22o_1
XU$$3399 U$$3399/A U$$3417/B VGND VGND VPWR VPWR U$$3399/X sky130_fd_sc_hd__xor2_1
XFILLER_34_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2654 U$$2654/A U$$2668/B VGND VGND VPWR VPWR U$$2654/X sky130_fd_sc_hd__xor2_1
XU$$2665 U$$2665/A1 U$$2665/A2 U$$2665/B1 U$$2665/B2 VGND VGND VPWR VPWR U$$2666/A
+ sky130_fd_sc_hd__a22o_1
XU$$1920 U$$2043/B VGND VGND VPWR VPWR U$$1920/Y sky130_fd_sc_hd__inv_1
XU$$1931 U$$1931/A U$$2007/B VGND VGND VPWR VPWR U$$1931/X sky130_fd_sc_hd__xor2_1
XU$$2676 U$$2676/A U$$2739/A VGND VGND VPWR VPWR U$$2676/X sky130_fd_sc_hd__xor2_1
XFILLER_34_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1942 U$$709/A1 U$$1986/A2 U$$709/B1 U$$1986/B2 VGND VGND VPWR VPWR U$$1943/A sky130_fd_sc_hd__a22o_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2687 U$$4331/A1 U$$2737/A2 U$$4196/A1 U$$2737/B2 VGND VGND VPWR VPWR U$$2688/A
+ sky130_fd_sc_hd__a22o_1
XU$$1953 U$$1953/A U$$1963/B VGND VGND VPWR VPWR U$$1953/X sky130_fd_sc_hd__xor2_1
XU$$2698 U$$2698/A U$$2708/B VGND VGND VPWR VPWR U$$2698/X sky130_fd_sc_hd__xor2_1
XU$$1964 U$$868/A1 U$$1964/A2 U$$868/B1 U$$1964/B2 VGND VGND VPWR VPWR U$$1965/A sky130_fd_sc_hd__a22o_1
XFILLER_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1975 U$$1975/A U$$1981/B VGND VGND VPWR VPWR U$$1975/X sky130_fd_sc_hd__xor2_1
XU$$1986 U$$616/A1 U$$1986/A2 U$$481/A1 U$$1986/B2 VGND VGND VPWR VPWR U$$1987/A sky130_fd_sc_hd__a22o_1
XFILLER_33_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1997 U$$1997/A U$$2031/B VGND VGND VPWR VPWR U$$1997/X sky130_fd_sc_hd__xor2_1
XFILLER_174_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_98_1 dadda_fa_5_98_1/A dadda_fa_5_98_1/B dadda_fa_5_98_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_99_0/B dadda_fa_7_98_0/A sky130_fd_sc_hd__fa_1
XFILLER_135_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$605 final_adder.U$$604/B final_adder.U$$489/X final_adder.U$$481/X
+ VGND VGND VPWR VPWR final_adder.U$$605/X sky130_fd_sc_hd__a21o_1
XFILLER_111_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$616 final_adder.U$$616/A final_adder.U$$616/B VGND VGND VPWR VPWR
+ final_adder.U$$720/A sky130_fd_sc_hd__and2_1
XFILLER_69_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$638 final_adder.U$$654/B final_adder.U$$638/B VGND VGND VPWR VPWR
+ final_adder.U$$750/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$649 final_adder.U$$648/B final_adder.U$$545/X final_adder.U$$529/X
+ VGND VGND VPWR VPWR final_adder.U$$649/X sky130_fd_sc_hd__a21o_1
XFILLER_57_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$60 U$$60/A1 U$$96/A2 U$$62/A1 U$$96/B2 VGND VGND VPWR VPWR U$$61/A sky130_fd_sc_hd__a22o_1
XU$$71 U$$71/A U$$87/B VGND VGND VPWR VPWR U$$71/X sky130_fd_sc_hd__xor2_1
XU$$82 U$$82/A1 U$$86/A2 U$$82/B1 U$$86/B2 VGND VGND VPWR VPWR U$$83/A sky130_fd_sc_hd__a22o_1
XU$$93 U$$93/A U$$97/B VGND VGND VPWR VPWR U$$93/X sky130_fd_sc_hd__xor2_1
XFILLER_25_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_93_0 dadda_fa_4_93_0/A dadda_fa_4_93_0/B dadda_fa_4_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_94_0/A dadda_fa_5_93_1/A sky130_fd_sc_hd__fa_1
XFILLER_153_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_107_2 U$$4211/X U$$4344/X U$$4477/X VGND VGND VPWR VPWR dadda_fa_4_108_1/A
+ dadda_fa_4_107_2/B sky130_fd_sc_hd__fa_1
XFILLER_137_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1205 U$$1205/A U$$1231/B VGND VGND VPWR VPWR U$$1205/X sky130_fd_sc_hd__xor2_1
XU$$1216 U$$120/A1 U$$1226/A2 U$$120/B1 U$$1226/B2 VGND VGND VPWR VPWR U$$1217/A sky130_fd_sc_hd__a22o_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1227 U$$1227/A U$$1227/B VGND VGND VPWR VPWR U$$1227/X sky130_fd_sc_hd__xor2_1
XU$$1238 U$$1236/B U$$1233/A input10/X U$$1233/Y VGND VGND VPWR VPWR U$$1238/X sky130_fd_sc_hd__a22o_1
XFILLER_43_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1249 U$$3030/A1 U$$1311/A2 U$$3030/B1 U$$1311/B2 VGND VGND VPWR VPWR U$$1250/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_102_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1021 final_adder.U$$4/SUM final_adder.U$$381/X final_adder.U$$4/COUT
+ VGND VGND VPWR VPWR final_adder.U$$1029/B sky130_fd_sc_hd__a21o_1
XFILLER_156_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1032 final_adder.U$$8/SUM final_adder.U$$503/X VGND VGND VPWR VPWR
+ output373/A sky130_fd_sc_hd__xor2_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1043 final_adder.U$$236/B final_adder.U$$1043/B VGND VGND VPWR VPWR
+ output295/A sky130_fd_sc_hd__xor2_1
XFILLER_144_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1054 final_adder.U$$224/A final_adder.U$$725/X VGND VGND VPWR VPWR
+ output308/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1065 final_adder.U$$214/B final_adder.U$$985/X VGND VGND VPWR VPWR
+ output320/A sky130_fd_sc_hd__xor2_1
XFILLER_109_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1076 final_adder.U$$202/A final_adder.U$$815/X VGND VGND VPWR VPWR
+ output332/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1087 final_adder.U$$192/B final_adder.U$$963/X VGND VGND VPWR VPWR
+ output344/A sky130_fd_sc_hd__xor2_1
XFILLER_109_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1098 final_adder.U$$180/A final_adder.U$$889/X VGND VGND VPWR VPWR
+ output356/A sky130_fd_sc_hd__xor2_1
XFILLER_124_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1350 U$$3391/B VGND VGND VPWR VPWR U$$3349/B sky130_fd_sc_hd__buf_8
XFILLER_39_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1361 U$$3287/A VGND VGND VPWR VPWR U$$3284/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_50_4 dadda_fa_2_50_4/A dadda_fa_2_50_4/B dadda_fa_2_50_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_1/CIN dadda_fa_3_50_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1372 U$$3123/B VGND VGND VPWR VPWR U$$3119/B sky130_fd_sc_hd__buf_4
Xfanout1383 fanout1391/X VGND VGND VPWR VPWR U$$2799/B sky130_fd_sc_hd__buf_6
Xfanout1394 U$$273/A VGND VGND VPWR VPWR U$$274/A sky130_fd_sc_hd__buf_4
XFILLER_66_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_43_3 dadda_fa_2_43_3/A dadda_fa_2_43_3/B dadda_fa_2_43_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_44_1/B dadda_fa_3_43_3/B sky130_fd_sc_hd__fa_1
XU$$3130 U$$3815/A1 U$$3144/A2 U$$3817/A1 U$$3144/B2 VGND VGND VPWR VPWR U$$3131/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3141 U$$3141/A U$$3147/B VGND VGND VPWR VPWR U$$3141/X sky130_fd_sc_hd__xor2_1
XU$$3152 input41/X VGND VGND VPWR VPWR U$$3154/B sky130_fd_sc_hd__inv_1
XU$$3163 U$$3163/A1 U$$3199/A2 U$$3163/B1 U$$3199/B2 VGND VGND VPWR VPWR U$$3164/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_36_2 U$$1542/X U$$1675/X U$$1808/X VGND VGND VPWR VPWR dadda_fa_3_37_1/A
+ dadda_fa_3_36_3/A sky130_fd_sc_hd__fa_1
XFILLER_46_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3174 U$$3174/A U$$3210/B VGND VGND VPWR VPWR U$$3174/X sky130_fd_sc_hd__xor2_1
XU$$2440 U$$2440/A U$$2466/A VGND VGND VPWR VPWR U$$2440/X sky130_fd_sc_hd__xor2_1
XU$$3185 U$$854/B1 U$$3207/A2 U$$721/A1 U$$3207/B2 VGND VGND VPWR VPWR U$$3186/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_13_1 dadda_fa_5_13_1/A dadda_fa_5_13_1/B dadda_ha_4_13_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_14_0/B dadda_fa_7_13_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_29_1 U$$464/X U$$597/X U$$730/X VGND VGND VPWR VPWR dadda_fa_3_30_1/CIN
+ dadda_fa_3_29_3/B sky130_fd_sc_hd__fa_1
XU$$3196 U$$3196/A U$$3196/B VGND VGND VPWR VPWR U$$3196/X sky130_fd_sc_hd__xor2_1
XU$$2451 U$$4367/B1 U$$2459/A2 U$$4234/A1 U$$2459/B2 VGND VGND VPWR VPWR U$$2452/A
+ sky130_fd_sc_hd__a22o_1
XU$$2462 U$$2462/A U$$2465/A VGND VGND VPWR VPWR U$$2462/X sky130_fd_sc_hd__xor2_1
XFILLER_50_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2473 U$$2473/A U$$2545/B VGND VGND VPWR VPWR U$$2473/X sky130_fd_sc_hd__xor2_1
XU$$2484 U$$2758/A1 U$$2532/A2 U$$2758/B1 U$$2532/B2 VGND VGND VPWR VPWR U$$2485/A
+ sky130_fd_sc_hd__a22o_1
XU$$2495 U$$2495/A U$$2529/B VGND VGND VPWR VPWR U$$2495/X sky130_fd_sc_hd__xor2_1
XU$$1750 U$$517/A1 U$$1758/A2 U$$517/B1 U$$1758/B2 VGND VGND VPWR VPWR U$$1751/A sky130_fd_sc_hd__a22o_1
XU$$1761 U$$1761/A U$$1761/B VGND VGND VPWR VPWR U$$1761/X sky130_fd_sc_hd__xor2_1
XFILLER_107_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1772 U$$2183/A1 U$$1778/A2 U$$4512/B1 U$$1778/B2 VGND VGND VPWR VPWR U$$1773/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1783 U$$1910/B VGND VGND VPWR VPWR U$$1783/Y sky130_fd_sc_hd__inv_1
XU$$1794 U$$1794/A U$$1828/B VGND VGND VPWR VPWR U$$1794/X sky130_fd_sc_hd__xor2_1
XFILLER_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput60 a[63] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput71 b[15] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput82 b[25] VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__buf_4
Xinput93 b[35] VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$402 final_adder.U$$406/B final_adder.U$$402/B VGND VGND VPWR VPWR
+ final_adder.U$$526/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$413 final_adder.U$$412/B final_adder.U$$291/X final_adder.U$$287/X
+ VGND VGND VPWR VPWR final_adder.U$$413/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$424 final_adder.U$$428/B final_adder.U$$424/B VGND VGND VPWR VPWR
+ final_adder.U$$548/B sky130_fd_sc_hd__and2_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$435 final_adder.U$$434/B final_adder.U$$313/X final_adder.U$$309/X
+ VGND VGND VPWR VPWR final_adder.U$$435/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$446 final_adder.U$$450/B final_adder.U$$446/B VGND VGND VPWR VPWR
+ final_adder.U$$570/B sky130_fd_sc_hd__and2_1
XFILLER_85_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$457 final_adder.U$$456/B final_adder.U$$335/X final_adder.U$$331/X
+ VGND VGND VPWR VPWR final_adder.U$$457/X sky130_fd_sc_hd__a21o_1
XFILLER_123_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$468 final_adder.U$$472/B final_adder.U$$468/B VGND VGND VPWR VPWR
+ final_adder.U$$592/B sky130_fd_sc_hd__and2_1
XU$$307 U$$307/A U$$339/B VGND VGND VPWR VPWR U$$307/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$479 final_adder.U$$478/B final_adder.U$$357/X final_adder.U$$353/X
+ VGND VGND VPWR VPWR final_adder.U$$479/X sky130_fd_sc_hd__a21o_1
XU$$318 U$$866/A1 U$$352/A2 U$$868/A1 U$$352/B2 VGND VGND VPWR VPWR U$$319/A sky130_fd_sc_hd__a22o_1
XU$$329 U$$329/A U$$363/B VGND VGND VPWR VPWR U$$329/X sky130_fd_sc_hd__xor2_1
XFILLER_38_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1012 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_112_0 dadda_fa_3_112_0/A U$$3423/X U$$3556/X VGND VGND VPWR VPWR dadda_fa_4_113_1/B
+ dadda_fa_4_112_2/A sky130_fd_sc_hd__fa_1
XFILLER_79_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_60_3 dadda_fa_3_60_3/A dadda_fa_3_60_3/B dadda_fa_3_60_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_1/B dadda_fa_4_60_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_53_2 dadda_fa_3_53_2/A dadda_fa_3_53_2/B dadda_fa_3_53_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_1/A dadda_fa_4_53_2/B sky130_fd_sc_hd__fa_1
XFILLER_0_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_69_2 U$$1209/X U$$1342/X U$$1475/X VGND VGND VPWR VPWR dadda_fa_1_70_6/CIN
+ dadda_fa_1_69_8/B sky130_fd_sc_hd__fa_1
XFILLER_75_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_46_1 dadda_fa_3_46_1/A dadda_fa_3_46_1/B dadda_fa_3_46_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_0/CIN dadda_fa_4_46_2/A sky130_fd_sc_hd__fa_1
XFILLER_76_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_23_0 dadda_fa_6_23_0/A dadda_fa_6_23_0/B dadda_fa_6_23_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_24_0/B dadda_fa_7_23_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_39_0 dadda_fa_3_39_0/A dadda_fa_3_39_0/B dadda_fa_3_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_0/B dadda_fa_4_39_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$991 final_adder.U$$220/A final_adder.U$$833/X final_adder.U$$991/B1
+ VGND VGND VPWR VPWR final_adder.U$$991/X sky130_fd_sc_hd__a21o_1
XU$$830 U$$8/A1 U$$876/A2 U$$8/B1 U$$876/B2 VGND VGND VPWR VPWR U$$831/A sky130_fd_sc_hd__a22o_1
XFILLER_63_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$841 U$$841/A U$$875/B VGND VGND VPWR VPWR U$$841/X sky130_fd_sc_hd__xor2_1
XU$$852 U$$987/B1 U$$904/A2 U$$852/B1 U$$904/B2 VGND VGND VPWR VPWR U$$853/A sky130_fd_sc_hd__a22o_1
XU$$863 U$$863/A U$$895/B VGND VGND VPWR VPWR U$$863/X sky130_fd_sc_hd__xor2_1
XU$$1002 U$$1002/A U$$982/B VGND VGND VPWR VPWR U$$1002/X sky130_fd_sc_hd__xor2_1
XU$$1013 U$$739/A1 U$$981/A2 U$$741/A1 U$$981/B2 VGND VGND VPWR VPWR U$$1014/A sky130_fd_sc_hd__a22o_1
XU$$874 U$$874/A1 U$$876/A2 U$$876/A1 U$$876/B2 VGND VGND VPWR VPWR U$$875/A sky130_fd_sc_hd__a22o_1
XU$$1024 U$$1024/A U$$998/B VGND VGND VPWR VPWR U$$1024/X sky130_fd_sc_hd__xor2_1
XFILLER_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$885 U$$885/A U$$925/B VGND VGND VPWR VPWR U$$885/X sky130_fd_sc_hd__xor2_1
XFILLER_17_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1035 U$$898/A1 U$$999/A2 U$$487/B1 U$$999/B2 VGND VGND VPWR VPWR U$$1036/A sky130_fd_sc_hd__a22o_1
XFILLER_90_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$896 U$$896/A1 U$$902/A2 U$$898/A1 U$$902/B2 VGND VGND VPWR VPWR U$$897/A sky130_fd_sc_hd__a22o_1
XU$$1046 U$$1046/A U$$1046/B VGND VGND VPWR VPWR U$$1046/X sky130_fd_sc_hd__xor2_1
XU$$1057 U$$98/A1 U$$997/A2 U$$98/B1 U$$997/B2 VGND VGND VPWR VPWR U$$1058/A sky130_fd_sc_hd__a22o_1
XFILLER_31_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_957 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1068 U$$1068/A U$$962/A VGND VGND VPWR VPWR U$$1068/X sky130_fd_sc_hd__xor2_1
XU$$1079 U$$120/A1 U$$1093/A2 U$$120/B1 U$$1093/B2 VGND VGND VPWR VPWR U$$1080/A sky130_fd_sc_hd__a22o_1
XFILLER_12_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_98_4 U$$3927/X U$$4060/X U$$4193/X VGND VGND VPWR VPWR dadda_fa_3_99_2/A
+ dadda_fa_3_98_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout609 U$$1758/A2 VGND VGND VPWR VPWR U$$1778/A2 sky130_fd_sc_hd__clkbuf_4
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1180 U$$4422/A1 VGND VGND VPWR VPWR U$$4420/B1 sky130_fd_sc_hd__buf_6
Xfanout1191 U$$4283/A1 VGND VGND VPWR VPWR U$$3048/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_54_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_41_0 U$$1552/X U$$1685/X U$$1818/X VGND VGND VPWR VPWR dadda_fa_3_42_0/B
+ dadda_fa_3_41_2/B sky130_fd_sc_hd__fa_1
XFILLER_23_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2270 U$$487/B1 U$$2272/A2 U$$902/A1 U$$2272/B2 VGND VGND VPWR VPWR U$$2271/A sky130_fd_sc_hd__a22o_1
XFILLER_50_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2281 U$$2281/A U$$2283/B VGND VGND VPWR VPWR U$$2281/X sky130_fd_sc_hd__xor2_1
XU$$2292 U$$2840/A1 U$$2310/A2 U$$2840/B1 U$$2310/B2 VGND VGND VPWR VPWR U$$2293/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1580 U$$1580/A U$$1584/B VGND VGND VPWR VPWR U$$1580/X sky130_fd_sc_hd__xor2_1
XFILLER_33_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1591 U$$632/A1 U$$1593/A2 U$$632/B1 U$$1593/B2 VGND VGND VPWR VPWR U$$1592/A sky130_fd_sc_hd__a22o_1
XFILLER_33_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_70_2 dadda_fa_4_70_2/A dadda_fa_4_70_2/B dadda_fa_4_70_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_71_0/CIN dadda_fa_5_70_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_86_2 U$$2307/X U$$2440/X U$$2573/X VGND VGND VPWR VPWR dadda_fa_2_87_3/B
+ dadda_fa_2_86_5/A sky130_fd_sc_hd__fa_1
XFILLER_143_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_63_1 dadda_fa_4_63_1/A dadda_fa_4_63_1/B dadda_fa_4_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_64_0/B dadda_fa_5_63_1/B sky130_fd_sc_hd__fa_1
XFILLER_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_79_1 U$$1495/X U$$1628/X U$$1761/X VGND VGND VPWR VPWR dadda_fa_2_80_0/CIN
+ dadda_fa_2_79_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_131_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_40_0 dadda_fa_7_40_0/A dadda_fa_7_40_0/B dadda_fa_7_40_0/CIN VGND VGND
+ VPWR VPWR _337_/D _208_/D sky130_fd_sc_hd__fa_1
XFILLER_103_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_56_0 dadda_fa_4_56_0/A dadda_fa_4_56_0/B dadda_fa_4_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_57_0/A dadda_fa_5_56_1/A sky130_fd_sc_hd__fa_1
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$210 final_adder.U$$210/A final_adder.U$$210/B VGND VGND VPWR VPWR
+ final_adder.U$$338/B sky130_fd_sc_hd__and2_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$221 final_adder.U$$220/B final_adder.U$$991/B1 final_adder.U$$221/B1
+ VGND VGND VPWR VPWR final_adder.U$$221/X sky130_fd_sc_hd__a21o_1
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$232 final_adder.U$$232/A final_adder.U$$232/B VGND VGND VPWR VPWR
+ final_adder.U$$360/B sky130_fd_sc_hd__and2_1
XFILLER_40_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$243 final_adder.U$$242/B final_adder.U$$243/A2 final_adder.U$$243/B1
+ VGND VGND VPWR VPWR final_adder.U$$243/X sky130_fd_sc_hd__a21o_1
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$265 final_adder.U$$264/B final_adder.U$$139/X final_adder.U$$137/X
+ VGND VGND VPWR VPWR final_adder.U$$265/X sky130_fd_sc_hd__a21o_1
XU$$104 U$$926/A1 U$$98/A2 U$$928/A1 U$$98/B2 VGND VGND VPWR VPWR U$$105/A sky130_fd_sc_hd__a22o_1
XFILLER_73_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$276 final_adder.U$$278/B final_adder.U$$276/B VGND VGND VPWR VPWR
+ final_adder.U$$402/B sky130_fd_sc_hd__and2_1
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$115 U$$115/A U$$121/B VGND VGND VPWR VPWR U$$115/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$287 final_adder.U$$286/B final_adder.U$$161/X final_adder.U$$159/X
+ VGND VGND VPWR VPWR final_adder.U$$287/X sky130_fd_sc_hd__a21o_1
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$126 U$$672/B1 U$$98/A2 U$$539/A1 U$$98/B2 VGND VGND VPWR VPWR U$$127/A sky130_fd_sc_hd__a22o_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$298 final_adder.U$$300/B final_adder.U$$298/B VGND VGND VPWR VPWR
+ final_adder.U$$424/B sky130_fd_sc_hd__and2_1
XFILLER_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$137 U$$3/A VGND VGND VPWR VPWR U$$137/Y sky130_fd_sc_hd__inv_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$148 U$$148/A U$$180/B VGND VGND VPWR VPWR U$$148/X sky130_fd_sc_hd__xor2_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$159 U$$22/A1 U$$213/A2 U$$24/A1 U$$213/B2 VGND VGND VPWR VPWR U$$160/A sky130_fd_sc_hd__a22o_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_392_ _397_/CLK _392_/D VGND VGND VPWR VPWR _392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_74_0 dadda_fa_0_74_0/A U$$820/X U$$953/X VGND VGND VPWR VPWR dadda_fa_1_75_7/CIN
+ dadda_fa_1_74_8/B sky130_fd_sc_hd__fa_1
XFILLER_49_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput250 c[94] VGND VGND VPWR VPWR input250/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$660 U$$934/A1 U$$674/A2 U$$936/A1 U$$674/B2 VGND VGND VPWR VPWR U$$661/A sky130_fd_sc_hd__a22o_1
XU$$671 U$$671/A U$$685/A VGND VGND VPWR VPWR U$$671/X sky130_fd_sc_hd__xor2_1
XFILLER_44_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$682 U$$956/A1 U$$682/A2 U$$682/B1 U$$682/B2 VGND VGND VPWR VPWR U$$683/A sky130_fd_sc_hd__a22o_1
XU$$693 U$$8/A1 U$$743/A2 U$$10/A1 U$$743/B2 VGND VGND VPWR VPWR U$$694/A sky130_fd_sc_hd__a22o_1
XFILLER_16_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_80_1 dadda_fa_5_80_1/A dadda_fa_5_80_1/B dadda_fa_5_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_81_0/B dadda_fa_7_80_0/A sky130_fd_sc_hd__fa_2
XFILLER_173_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_96_1 U$$2859/X U$$2992/X U$$3125/X VGND VGND VPWR VPWR dadda_fa_3_97_0/CIN
+ dadda_fa_3_96_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_73_0 dadda_fa_5_73_0/A dadda_fa_5_73_0/B dadda_fa_5_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_74_0/A dadda_fa_6_73_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_126_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_98_0_1935 VGND VGND VPWR VPWR dadda_fa_2_98_0/A dadda_fa_2_98_0_1935/LO
+ sky130_fd_sc_hd__conb_1
Xdadda_fa_2_89_0 U$$3377/X U$$3510/X U$$3643/X VGND VGND VPWR VPWR dadda_fa_3_90_0/B
+ dadda_fa_3_89_2/B sky130_fd_sc_hd__fa_1
XFILLER_99_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout406 U$$819/A2 VGND VGND VPWR VPWR U$$817/A2 sky130_fd_sc_hd__buf_6
Xfanout417 U$$4309/A2 VGND VGND VPWR VPWR U$$4289/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout428 U$$415/X VGND VGND VPWR VPWR U$$543/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_72_8 dadda_fa_1_72_8/A dadda_fa_1_72_8/B dadda_fa_1_72_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_73_3/A dadda_fa_3_72_0/A sky130_fd_sc_hd__fa_2
XFILLER_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout439 U$$4190/A2 VGND VGND VPWR VPWR U$$4226/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_140_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_65_7 dadda_fa_1_65_7/A dadda_fa_1_65_7/B dadda_fa_1_65_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_66_2/CIN dadda_fa_2_65_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_58_6 U$$3980/X U$$4006/B input210/X VGND VGND VPWR VPWR dadda_fa_2_59_2/B
+ dadda_fa_2_58_5/B sky130_fd_sc_hd__fa_1
XFILLER_100_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_1_92_2 U$$2718/X U$$2851/X VGND VGND VPWR VPWR dadda_fa_2_93_5/B dadda_fa_3_92_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_109_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_88_0 dadda_fa_7_88_0/A dadda_fa_7_88_0/B dadda_fa_7_88_0/CIN VGND VGND
+ VPWR VPWR _385_/D _256_/D sky130_fd_sc_hd__fa_1
XFILLER_89_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_91_0 U$$1917/Y U$$2051/X U$$2184/X VGND VGND VPWR VPWR dadda_fa_2_92_4/B
+ dadda_fa_2_91_5/B sky130_fd_sc_hd__fa_1
XFILLER_135_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout940 U$$2480/A1 VGND VGND VPWR VPWR U$$3163/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout951 fanout957/X VGND VGND VPWR VPWR U$$3372/B1 sky130_fd_sc_hd__buf_4
XU$$4408 U$$4408/A1 U$$4388/X U$$4410/A1 U$$4458/B2 VGND VGND VPWR VPWR U$$4409/A
+ sky130_fd_sc_hd__a22o_1
Xfanout962 fanout966/X VGND VGND VPWR VPWR U$$82/B1 sky130_fd_sc_hd__buf_6
XU$$4419 U$$4419/A U$$4419/B VGND VGND VPWR VPWR U$$4419/X sky130_fd_sc_hd__xor2_1
Xfanout973 U$$4466/A1 VGND VGND VPWR VPWR U$$4464/B1 sky130_fd_sc_hd__buf_4
Xfanout984 input94/X VGND VGND VPWR VPWR fanout984/X sky130_fd_sc_hd__buf_8
Xfanout995 fanout999/A VGND VGND VPWR VPWR U$$487/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3707 U$$3979/B1 U$$3703/X U$$3846/A1 U$$3704/X VGND VGND VPWR VPWR U$$3708/A sky130_fd_sc_hd__a22o_1
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3718 U$$3718/A U$$3734/B VGND VGND VPWR VPWR U$$3718/X sky130_fd_sc_hd__xor2_1
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3729 U$$4001/B1 U$$3757/A2 U$$854/A1 U$$3757/B2 VGND VGND VPWR VPWR U$$3730/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_103_0 dadda_fa_6_103_0/A dadda_fa_6_103_0/B dadda_fa_6_103_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_104_0/B dadda_fa_7_103_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_23_3 U$$1516/X input172/X dadda_fa_3_23_3/CIN VGND VGND VPWR VPWR dadda_fa_4_24_1/B
+ dadda_fa_4_23_2/CIN sky130_fd_sc_hd__fa_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_375_ _375_/CLK _375_/D VGND VGND VPWR VPWR _375_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_90_0 dadda_fa_6_90_0/A dadda_fa_6_90_0/B dadda_fa_6_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_91_0/B dadda_fa_7_90_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_70_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_68_5 dadda_fa_2_68_5/A dadda_fa_2_68_5/B dadda_fa_2_68_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_2/A dadda_fa_4_68_0/A sky130_fd_sc_hd__fa_1
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$490 U$$490/A U$$498/B VGND VGND VPWR VPWR U$$490/X sky130_fd_sc_hd__xor2_1
XFILLER_149_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2198_1800 VGND VGND VPWR VPWR U$$2198_1800/HI U$$2198/A1 sky130_fd_sc_hd__conb_1
XFILLER_160_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_70_5 U$$4270/X U$$4403/X input224/X VGND VGND VPWR VPWR dadda_fa_2_71_2/A
+ dadda_fa_2_70_5/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_63_4 U$$3990/X U$$4123/X U$$4256/X VGND VGND VPWR VPWR dadda_fa_2_64_1/CIN
+ dadda_fa_2_63_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_75_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_56_3 U$$2380/X U$$2513/X U$$2646/X VGND VGND VPWR VPWR dadda_fa_2_57_1/B
+ dadda_fa_2_56_4/B sky130_fd_sc_hd__fa_1
Xdadda_fa_4_33_2 dadda_fa_4_33_2/A dadda_fa_4_33_2/B dadda_fa_4_33_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_34_0/CIN dadda_fa_5_33_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_49_2 U$$903/X U$$1036/X U$$1169/X VGND VGND VPWR VPWR dadda_fa_2_50_1/B
+ dadda_fa_2_49_4/B sky130_fd_sc_hd__fa_1
XFILLER_82_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_26_1 dadda_fa_4_26_1/A dadda_fa_4_26_1/B dadda_fa_4_26_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_27_0/B dadda_fa_5_26_1/B sky130_fd_sc_hd__fa_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_19_0 U$$1109/X U$$1242/X input167/X VGND VGND VPWR VPWR dadda_fa_5_20_0/A
+ dadda_fa_5_19_1/A sky130_fd_sc_hd__fa_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1702 U$$2844/B1 VGND VGND VPWR VPWR U$$928/A1 sky130_fd_sc_hd__buf_6
XFILLER_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1713 fanout1718/X VGND VGND VPWR VPWR U$$787/B1 sky130_fd_sc_hd__buf_6
Xfanout1724 U$$4486/A1 VGND VGND VPWR VPWR U$$4349/A1 sky130_fd_sc_hd__buf_4
Xfanout1735 U$$370/B1 VGND VGND VPWR VPWR U$$98/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1746 U$$505/B1 VGND VGND VPWR VPWR U$$3110/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1757 U$$914/B1 VGND VGND VPWR VPWR U$$916/A1 sky130_fd_sc_hd__buf_6
XU$$4205 U$$4205/A U$$4227/B VGND VGND VPWR VPWR U$$4205/X sky130_fd_sc_hd__xor2_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout770 U$$3072/B2 VGND VGND VPWR VPWR U$$3066/B2 sky130_fd_sc_hd__buf_4
XU$$4216 U$$4353/A1 U$$4240/A2 U$$4353/B1 U$$4240/B2 VGND VGND VPWR VPWR U$$4217/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1768 U$$3515/B1 VGND VGND VPWR VPWR U$$4474/B1 sky130_fd_sc_hd__buf_2
Xfanout781 U$$2977/B2 VGND VGND VPWR VPWR U$$2979/B2 sky130_fd_sc_hd__buf_4
XU$$4227 U$$4227/A U$$4227/B VGND VGND VPWR VPWR U$$4227/X sky130_fd_sc_hd__xor2_1
Xfanout1779 input100/X VGND VGND VPWR VPWR U$$912/A1 sky130_fd_sc_hd__buf_4
XFILLER_59_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4238 U$$4375/A1 U$$4240/A2 U$$4375/B1 U$$4240/B2 VGND VGND VPWR VPWR U$$4239/A
+ sky130_fd_sc_hd__a22o_1
Xfanout792 U$$346/B2 VGND VGND VPWR VPWR U$$340/B2 sky130_fd_sc_hd__buf_2
XU$$3504 U$$3504/A U$$3506/B VGND VGND VPWR VPWR U$$3504/X sky130_fd_sc_hd__xor2_1
XFILLER_65_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4249 U$$4383/A VGND VGND VPWR VPWR U$$4249/Y sky130_fd_sc_hd__inv_1
XFILLER_92_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3515 U$$3650/B1 U$$3557/A2 U$$3515/B1 U$$3557/B2 VGND VGND VPWR VPWR U$$3516/A
+ sky130_fd_sc_hd__a22o_1
XU$$3526 U$$3526/A U$$3548/B VGND VGND VPWR VPWR U$$3526/X sky130_fd_sc_hd__xor2_1
XFILLER_74_941 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3537 U$$4359/A1 U$$3549/A2 U$$3948/B1 U$$3549/B2 VGND VGND VPWR VPWR U$$3538/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2803 U$$2803/A U$$2877/A VGND VGND VPWR VPWR U$$2803/X sky130_fd_sc_hd__xor2_1
XU$$3548 U$$3548/A U$$3548/B VGND VGND VPWR VPWR U$$3548/X sky130_fd_sc_hd__xor2_1
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3559 U$$3559/A1 U$$3559/A2 U$$3559/B1 U$$3559/B2 VGND VGND VPWR VPWR U$$3560/A
+ sky130_fd_sc_hd__a22o_1
XU$$2814 U$$2814/A1 U$$2856/A2 U$$74/B1 U$$2856/B2 VGND VGND VPWR VPWR U$$2815/A sky130_fd_sc_hd__a22o_1
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2825 U$$2825/A U$$2877/A VGND VGND VPWR VPWR U$$2825/X sky130_fd_sc_hd__xor2_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2836 U$$2973/A1 U$$2840/A2 U$$2973/B1 U$$2840/B2 VGND VGND VPWR VPWR U$$2837/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2847 U$$2847/A U$$2876/A VGND VGND VPWR VPWR U$$2847/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_21_0 U$$49/X U$$182/X U$$315/X VGND VGND VPWR VPWR dadda_fa_4_22_0/B dadda_fa_4_21_1/CIN
+ sky130_fd_sc_hd__fa_1
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2858 U$$2993/B1 U$$2872/A2 U$$2860/A1 U$$2872/B2 VGND VGND VPWR VPWR U$$2859/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2869 U$$2869/A U$$2871/B VGND VGND VPWR VPWR U$$2869/X sky130_fd_sc_hd__xor2_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_358_ _358_/CLK _358_/D VGND VGND VPWR VPWR _358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_289_ _420_/CLK _289_/D VGND VGND VPWR VPWR _289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_80_4 dadda_fa_2_80_4/A dadda_fa_2_80_4/B dadda_fa_2_80_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_1/CIN dadda_fa_3_80_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_73_3 dadda_fa_2_73_3/A dadda_fa_2_73_3/B dadda_fa_2_73_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_1/B dadda_fa_3_73_3/B sky130_fd_sc_hd__fa_1
XFILLER_123_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_66_2 dadda_fa_2_66_2/A dadda_fa_2_66_2/B dadda_fa_2_66_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_1/A dadda_fa_3_66_3/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$809 final_adder.U$$776/A final_adder.U$$729/X final_adder.U$$697/X
+ VGND VGND VPWR VPWR final_adder.U$$809/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_5_43_1 dadda_fa_5_43_1/A dadda_fa_5_43_1/B dadda_fa_5_43_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_44_0/B dadda_fa_7_43_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_59_1 dadda_fa_2_59_1/A dadda_fa_2_59_1/B dadda_fa_2_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_0/CIN dadda_fa_3_59_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_84_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 a[11] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_36_0 dadda_fa_5_36_0/A dadda_fa_5_36_0/B dadda_fa_5_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_37_0/A dadda_fa_6_36_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_149_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_110_0 dadda_fa_5_110_0/A dadda_fa_5_110_0/B dadda_fa_5_110_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_111_0/A dadda_fa_6_110_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$1 _297_/Q _169_/Q VGND VGND VPWR VPWR final_adder.U$$255/B1 final_adder.U$$1/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_69_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput340 output340/A VGND VGND VPWR VPWR o[5] sky130_fd_sc_hd__buf_2
XFILLER_134_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput351 output351/A VGND VGND VPWR VPWR o[6] sky130_fd_sc_hd__buf_2
Xoutput362 output362/A VGND VGND VPWR VPWR o[7] sky130_fd_sc_hd__buf_2
Xoutput373 output373/A VGND VGND VPWR VPWR o[8] sky130_fd_sc_hd__buf_2
Xoutput384 output384/A VGND VGND VPWR VPWR o[9] sky130_fd_sc_hd__buf_2
Xfanout1009 U$$4458/A1 VGND VGND VPWR VPWR U$$4456/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_160_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_61_1 U$$2390/X U$$2523/X U$$2656/X VGND VGND VPWR VPWR dadda_fa_2_62_0/CIN
+ dadda_fa_2_61_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_101_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_0 U$$780/X U$$913/X U$$1046/X VGND VGND VPWR VPWR dadda_fa_2_55_0/B
+ dadda_fa_2_54_3/B sky130_fd_sc_hd__fa_1
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1409 U$$1409/A U$$1449/B VGND VGND VPWR VPWR U$$1409/X sky130_fd_sc_hd__xor2_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_212_ _342_/CLK _212_/D VGND VGND VPWR VPWR _212_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_129_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_90_3 dadda_fa_3_90_3/A dadda_fa_3_90_3/B dadda_fa_3_90_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_1/B dadda_fa_4_90_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_136_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4515_1905 VGND VGND VPWR VPWR U$$4515_1905/HI U$$4515/B sky130_fd_sc_hd__conb_1
XFILLER_125_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_83_2 dadda_fa_3_83_2/A dadda_fa_3_83_2/B dadda_fa_3_83_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_1/A dadda_fa_4_83_2/B sky130_fd_sc_hd__fa_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_76_1 dadda_fa_3_76_1/A dadda_fa_3_76_1/B dadda_fa_3_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_0/CIN dadda_fa_4_76_2/A sky130_fd_sc_hd__fa_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_53_0 dadda_fa_6_53_0/A dadda_fa_6_53_0/B dadda_fa_6_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_54_0/B dadda_fa_7_53_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_69_0 dadda_fa_3_69_0/A dadda_fa_3_69_0/B dadda_fa_3_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_0/B dadda_fa_4_69_1/CIN sky130_fd_sc_hd__fa_1
Xfanout1510 U$$3314/A1 VGND VGND VPWR VPWR U$$709/B1 sky130_fd_sc_hd__buf_4
Xfanout1521 U$$4408/A1 VGND VGND VPWR VPWR U$$3447/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1532 U$$4404/A1 VGND VGND VPWR VPWR U$$2897/A1 sky130_fd_sc_hd__buf_4
Xfanout1543 U$$3833/A1 VGND VGND VPWR VPWR U$$4107/A1 sky130_fd_sc_hd__buf_4
Xfanout1554 input123/X VGND VGND VPWR VPWR U$$3692/B1 sky130_fd_sc_hd__buf_2
XU$$4002 U$$4002/A U$$4006/B VGND VGND VPWR VPWR U$$4002/X sky130_fd_sc_hd__xor2_1
Xfanout1565 U$$4512/A1 VGND VGND VPWR VPWR U$$539/A1 sky130_fd_sc_hd__buf_6
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4013 U$$4150/A1 U$$4057/A2 U$$4152/A1 U$$4057/B2 VGND VGND VPWR VPWR U$$4014/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4024 U$$4024/A U$$4040/B VGND VGND VPWR VPWR U$$4024/X sky130_fd_sc_hd__xor2_1
Xfanout1576 U$$4402/A1 VGND VGND VPWR VPWR U$$4400/B1 sky130_fd_sc_hd__buf_4
XU$$4035 U$$4307/B1 U$$4045/A2 U$$4174/A1 U$$4045/B2 VGND VGND VPWR VPWR U$$4036/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1587 U$$49/B VGND VGND VPWR VPWR U$$9/B sky130_fd_sc_hd__buf_4
Xfanout1598 U$$2729/A1 VGND VGND VPWR VPWR U$$3551/A1 sky130_fd_sc_hd__buf_4
XFILLER_65_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3301 U$$3301/A U$$3341/B VGND VGND VPWR VPWR U$$3301/X sky130_fd_sc_hd__xor2_1
XU$$4046 U$$4046/A U$$4110/A VGND VGND VPWR VPWR U$$4046/X sky130_fd_sc_hd__xor2_1
XFILLER_19_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3312 U$$4408/A1 U$$3390/A2 U$$4410/A1 U$$3390/B2 VGND VGND VPWR VPWR U$$3313/A
+ sky130_fd_sc_hd__a22o_1
XU$$4057 U$$4331/A1 U$$4057/A2 U$$4196/A1 U$$4057/B2 VGND VGND VPWR VPWR U$$4058/A
+ sky130_fd_sc_hd__a22o_1
XU$$4068 U$$4068/A U$$4094/B VGND VGND VPWR VPWR U$$4068/X sky130_fd_sc_hd__xor2_1
XU$$3323 U$$3323/A U$$3335/B VGND VGND VPWR VPWR U$$3323/X sky130_fd_sc_hd__xor2_1
XFILLER_93_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_112_2 dadda_fa_4_112_2/A dadda_fa_4_112_2/B dadda_ha_3_112_2/SUM VGND
+ VGND VPWR VPWR dadda_fa_5_113_0/CIN dadda_fa_5_112_1/CIN sky130_fd_sc_hd__fa_1
XU$$3334 U$$4430/A1 U$$3340/A2 U$$4158/A1 U$$3340/B2 VGND VGND VPWR VPWR U$$3335/A
+ sky130_fd_sc_hd__a22o_1
XU$$4079 U$$4214/B1 U$$4081/A2 U$$4081/A1 U$$4081/B2 VGND VGND VPWR VPWR U$$4080/A
+ sky130_fd_sc_hd__a22o_1
XU$$2600 U$$3285/A1 U$$2600/A2 U$$2600/B1 U$$2600/B2 VGND VGND VPWR VPWR U$$2601/A
+ sky130_fd_sc_hd__a22o_1
XU$$3345 U$$3345/A U$$3349/B VGND VGND VPWR VPWR U$$3345/X sky130_fd_sc_hd__xor2_1
XU$$3356 U$$3628/B1 U$$3372/A2 U$$3630/B1 U$$3372/B2 VGND VGND VPWR VPWR U$$3357/A
+ sky130_fd_sc_hd__a22o_1
XU$$2611 U$$2748/A1 U$$2681/A2 U$$3296/B1 U$$2681/B2 VGND VGND VPWR VPWR U$$2612/A
+ sky130_fd_sc_hd__a22o_1
XU$$2622 U$$2622/A U$$2662/B VGND VGND VPWR VPWR U$$2622/X sky130_fd_sc_hd__xor2_1
XU$$3367 U$$3367/A U$$3373/B VGND VGND VPWR VPWR U$$3367/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_105_1 dadda_fa_4_105_1/A dadda_fa_4_105_1/B dadda_fa_4_105_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_106_0/B dadda_fa_5_105_1/B sky130_fd_sc_hd__fa_1
XFILLER_18_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3378 U$$3650/B1 U$$3378/A2 U$$3515/B1 U$$3378/B2 VGND VGND VPWR VPWR U$$3379/A
+ sky130_fd_sc_hd__a22o_1
XU$$2633 U$$576/B1 U$$2681/A2 U$$443/A1 U$$2681/B2 VGND VGND VPWR VPWR U$$2634/A sky130_fd_sc_hd__a22o_1
XU$$2644 U$$2644/A U$$2724/B VGND VGND VPWR VPWR U$$2644/X sky130_fd_sc_hd__xor2_1
XU$$1910 U$$1910/A U$$1910/B VGND VGND VPWR VPWR U$$1910/X sky130_fd_sc_hd__xor2_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3389 U$$3389/A U$$3391/B VGND VGND VPWR VPWR U$$3389/X sky130_fd_sc_hd__xor2_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2655 U$$735/B1 U$$2665/A2 U$$602/A1 U$$2665/B2 VGND VGND VPWR VPWR U$$2656/A sky130_fd_sc_hd__a22o_1
XFILLER_34_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2666 U$$2666/A U$$2668/B VGND VGND VPWR VPWR U$$2666/X sky130_fd_sc_hd__xor2_1
XU$$1921 U$$2043/B U$$1921/B VGND VGND VPWR VPWR U$$1921/X sky130_fd_sc_hd__and2_1
XFILLER_92_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1932 U$$2480/A1 U$$1986/A2 U$$3030/A1 U$$1986/B2 VGND VGND VPWR VPWR U$$1933/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2677 U$$4456/B1 U$$2681/A2 U$$4049/A1 U$$2681/B2 VGND VGND VPWR VPWR U$$2678/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1943 U$$1943/A U$$1971/B VGND VGND VPWR VPWR U$$1943/X sky130_fd_sc_hd__xor2_1
XU$$2688 U$$2688/A U$$2738/B VGND VGND VPWR VPWR U$$2688/X sky130_fd_sc_hd__xor2_1
XU$$1954 U$$995/A1 U$$1964/A2 U$$997/A1 U$$1964/B2 VGND VGND VPWR VPWR U$$1955/A sky130_fd_sc_hd__a22o_1
XU$$2699 U$$2973/A1 U$$2707/A2 U$$2973/B1 U$$2707/B2 VGND VGND VPWR VPWR U$$2700/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1965 U$$1965/A U$$2007/B VGND VGND VPWR VPWR U$$1965/X sky130_fd_sc_hd__xor2_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1976 U$$878/B1 U$$1986/A2 U$$745/A1 U$$1986/B2 VGND VGND VPWR VPWR U$$1977/A sky130_fd_sc_hd__a22o_1
XU$$1987 U$$1987/A U$$2015/B VGND VGND VPWR VPWR U$$1987/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_126_0 dadda_fa_7_126_0/A dadda_fa_7_126_0/B dadda_fa_7_126_0/CIN VGND
+ VGND VPWR VPWR _423_/D _294_/D sky130_fd_sc_hd__fa_1
XU$$1998 U$$3503/B1 U$$2046/A2 U$$3370/A1 U$$2046/B2 VGND VGND VPWR VPWR U$$1999/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_71_0 dadda_fa_2_71_0/A dadda_fa_2_71_0/B dadda_fa_2_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_0/B dadda_fa_3_71_2/B sky130_fd_sc_hd__fa_1
XFILLER_97_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$606 final_adder.U$$614/B final_adder.U$$606/B VGND VGND VPWR VPWR
+ final_adder.U$$710/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$617 final_adder.U$$616/B final_adder.U$$501/X final_adder.U$$493/X
+ VGND VGND VPWR VPWR final_adder.U$$617/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$628 final_adder.U$$644/B final_adder.U$$628/B VGND VGND VPWR VPWR
+ final_adder.U$$740/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$639 final_adder.U$$638/B final_adder.U$$535/X final_adder.U$$519/X
+ VGND VGND VPWR VPWR final_adder.U$$639/X sky130_fd_sc_hd__a21o_1
XFILLER_72_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$50 U$$50/A1 U$$86/A2 U$$50/B1 U$$86/B2 VGND VGND VPWR VPWR U$$51/A sky130_fd_sc_hd__a22o_1
XU$$61 U$$61/A U$$97/B VGND VGND VPWR VPWR U$$61/X sky130_fd_sc_hd__xor2_1
XFILLER_53_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$72 U$$72/A1 U$$74/A2 U$$74/A1 U$$74/B2 VGND VGND VPWR VPWR U$$73/A sky130_fd_sc_hd__a22o_1
XFILLER_37_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$83 U$$83/A U$$87/B VGND VGND VPWR VPWR U$$83/X sky130_fd_sc_hd__xor2_1
XU$$94 U$$94/A1 U$$96/A2 U$$96/A1 U$$96/B2 VGND VGND VPWR VPWR U$$95/A sky130_fd_sc_hd__a22o_1
XFILLER_72_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3890 U$$4438/A1 U$$3906/A2 U$$4027/B1 U$$3906/B2 VGND VGND VPWR VPWR U$$3891/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_93_1 dadda_fa_4_93_1/A dadda_fa_4_93_1/B dadda_fa_4_93_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_94_0/B dadda_fa_5_93_1/B sky130_fd_sc_hd__fa_1
XFILLER_165_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_70_0 dadda_fa_7_70_0/A dadda_fa_7_70_0/B dadda_fa_7_70_0/CIN VGND VGND
+ VPWR VPWR _367_/D _238_/D sky130_fd_sc_hd__fa_1
XFILLER_118_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_86_0 dadda_fa_4_86_0/A dadda_fa_4_86_0/B dadda_fa_4_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_87_0/A dadda_fa_5_86_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_107_3 input137/X dadda_fa_3_107_3/B dadda_fa_3_107_3/CIN VGND VGND VPWR
+ VPWR dadda_fa_4_108_1/B dadda_fa_4_107_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$271_1807 VGND VGND VPWR VPWR U$$271_1807/HI U$$271/B1 sky130_fd_sc_hd__conb_1
XFILLER_43_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1206 U$$932/A1 U$$1230/A2 U$$934/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1207/A sky130_fd_sc_hd__a22o_1
XU$$1217 U$$1217/A U$$1227/B VGND VGND VPWR VPWR U$$1217/X sky130_fd_sc_hd__xor2_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1228 U$$678/B1 U$$1230/A2 U$$406/B1 U$$1230/B2 VGND VGND VPWR VPWR U$$1229/A sky130_fd_sc_hd__a22o_1
XU$$1239 U$$1239/A1 U$$1309/A2 U$$967/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1240/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1011 final_adder.U$$240/A final_adder.U$$621/X final_adder.U$$241/A2
+ VGND VGND VPWR VPWR final_adder.U$$1039/B sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$1033 final_adder.U$$9/SUM final_adder.U$$1033/B VGND VGND VPWR VPWR
+ output384/A sky130_fd_sc_hd__xor2_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1044 final_adder.U$$234/A final_adder.U$$735/X VGND VGND VPWR VPWR
+ output297/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1055 final_adder.U$$224/B final_adder.U$$995/X VGND VGND VPWR VPWR
+ output309/A sky130_fd_sc_hd__xor2_1
XFILLER_109_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1066 final_adder.U$$212/A final_adder.U$$825/X VGND VGND VPWR VPWR
+ output321/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1077 final_adder.U$$202/B final_adder.U$$973/X VGND VGND VPWR VPWR
+ output333/A sky130_fd_sc_hd__xor2_1
XFILLER_137_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1088 final_adder.U$$190/A final_adder.U$$803/X VGND VGND VPWR VPWR
+ output345/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1099 final_adder.U$$180/B final_adder.U$$951/X VGND VGND VPWR VPWR
+ output357/A sky130_fd_sc_hd__xor2_1
XFILLER_124_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1340 input47/X VGND VGND VPWR VPWR U$$3562/A sky130_fd_sc_hd__buf_6
XFILLER_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1351 U$$3424/A VGND VGND VPWR VPWR U$$3417/B sky130_fd_sc_hd__buf_6
XFILLER_38_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1362 U$$3287/A VGND VGND VPWR VPWR U$$3286/B sky130_fd_sc_hd__clkbuf_4
XFILLER_39_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_50_5 dadda_fa_2_50_5/A dadda_fa_2_50_5/B dadda_fa_2_50_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_2/A dadda_fa_4_50_0/A sky130_fd_sc_hd__fa_2
Xfanout1373 input40/X VGND VGND VPWR VPWR U$$3123/B sky130_fd_sc_hd__buf_6
Xfanout1384 fanout1391/X VGND VGND VPWR VPWR U$$2805/B sky130_fd_sc_hd__buf_6
XFILLER_93_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1395 U$$260/B VGND VGND VPWR VPWR U$$273/A sky130_fd_sc_hd__buf_4
Xdadda_fa_2_43_4 dadda_fa_2_43_4/A dadda_fa_2_43_4/B dadda_fa_2_43_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_44_1/CIN dadda_fa_3_43_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3120 U$$4214/B1 U$$3148/A2 U$$4081/A1 U$$3148/B2 VGND VGND VPWR VPWR U$$3121/A
+ sky130_fd_sc_hd__a22o_1
XU$$3131 U$$3131/A U$$3150/A VGND VGND VPWR VPWR U$$3131/X sky130_fd_sc_hd__xor2_1
XFILLER_47_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3142 U$$3416/A1 U$$3144/A2 U$$3418/A1 U$$3144/B2 VGND VGND VPWR VPWR U$$3143/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_ha_6_2_0 U$$11/X U$$144/X VGND VGND VPWR VPWR dadda_fa_7_3_0/B dadda_ha_6_2_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$3153 U$$3288/A VGND VGND VPWR VPWR U$$3153/Y sky130_fd_sc_hd__inv_1
XFILLER_35_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_36_3 U$$1941/X U$$2074/X U$$2207/X VGND VGND VPWR VPWR dadda_fa_3_37_1/B
+ dadda_fa_3_36_3/B sky130_fd_sc_hd__fa_1
XU$$3164 U$$3164/A U$$3196/B VGND VGND VPWR VPWR U$$3164/X sky130_fd_sc_hd__xor2_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2430 U$$2430/A U$$2466/A VGND VGND VPWR VPWR U$$2430/X sky130_fd_sc_hd__xor2_1
XU$$3175 U$$4408/A1 U$$3255/A2 U$$4410/A1 U$$3255/B2 VGND VGND VPWR VPWR U$$3176/A
+ sky130_fd_sc_hd__a22o_1
XU$$2441 U$$2576/B1 U$$2443/A2 U$$2578/B1 U$$2443/B2 VGND VGND VPWR VPWR U$$2442/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3186 U$$3186/A U$$3208/B VGND VGND VPWR VPWR U$$3186/X sky130_fd_sc_hd__xor2_1
XU$$3197 U$$4430/A1 U$$3207/A2 U$$4158/A1 U$$3207/B2 VGND VGND VPWR VPWR U$$3198/A
+ sky130_fd_sc_hd__a22o_1
XU$$2452 U$$2452/A U$$2456/B VGND VGND VPWR VPWR U$$2452/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_29_2 U$$863/X U$$996/X U$$1129/X VGND VGND VPWR VPWR dadda_fa_3_30_2/A
+ dadda_fa_3_29_3/CIN sky130_fd_sc_hd__fa_1
XU$$2463 input124/X U$$2463/A2 U$$2463/B1 U$$2463/B2 VGND VGND VPWR VPWR U$$2464/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2474 U$$967/A1 U$$2546/A2 U$$969/A1 U$$2546/B2 VGND VGND VPWR VPWR U$$2475/A sky130_fd_sc_hd__a22o_1
XU$$2485 U$$2485/A U$$2529/B VGND VGND VPWR VPWR U$$2485/X sky130_fd_sc_hd__xor2_1
XFILLER_61_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1740 U$$505/B1 U$$1774/A2 U$$370/B1 U$$1774/B2 VGND VGND VPWR VPWR U$$1741/A sky130_fd_sc_hd__a22o_1
XU$$2496 U$$2631/B1 U$$2540/A2 U$$852/B1 U$$2540/B2 VGND VGND VPWR VPWR U$$2497/A
+ sky130_fd_sc_hd__a22o_1
XU$$1751 U$$1751/A U$$1761/B VGND VGND VPWR VPWR U$$1751/X sky130_fd_sc_hd__xor2_1
XU$$1762 U$$2310/A1 U$$1778/A2 U$$942/A1 U$$1778/B2 VGND VGND VPWR VPWR U$$1763/A
+ sky130_fd_sc_hd__a22o_1
XU$$1773 U$$1773/A U$$1777/B VGND VGND VPWR VPWR U$$1773/X sky130_fd_sc_hd__xor2_1
XU$$1784 U$$1910/B U$$1784/B VGND VGND VPWR VPWR U$$1784/X sky130_fd_sc_hd__and2_1
XU$$1795 U$$2754/A1 U$$1831/A2 U$$2891/B1 U$$1831/B2 VGND VGND VPWR VPWR U$$1796/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput50 a[54] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput61 a[6] VGND VGND VPWR VPWR U$$412/A sky130_fd_sc_hd__buf_2
Xinput72 b[16] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput83 b[26] VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_4
Xinput94 b[36] VGND VGND VPWR VPWR input94/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$403 final_adder.U$$402/B final_adder.U$$281/X final_adder.U$$277/X
+ VGND VGND VPWR VPWR final_adder.U$$403/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$414 final_adder.U$$418/B final_adder.U$$414/B VGND VGND VPWR VPWR
+ final_adder.U$$538/B sky130_fd_sc_hd__and2_1
XFILLER_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$425 final_adder.U$$424/B final_adder.U$$303/X final_adder.U$$299/X
+ VGND VGND VPWR VPWR final_adder.U$$425/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$436 final_adder.U$$440/B final_adder.U$$436/B VGND VGND VPWR VPWR
+ final_adder.U$$560/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$447 final_adder.U$$446/B final_adder.U$$325/X final_adder.U$$321/X
+ VGND VGND VPWR VPWR final_adder.U$$447/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$458 final_adder.U$$462/B final_adder.U$$458/B VGND VGND VPWR VPWR
+ final_adder.U$$582/B sky130_fd_sc_hd__and2_1
XFILLER_85_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$469 final_adder.U$$468/B final_adder.U$$347/X final_adder.U$$343/X
+ VGND VGND VPWR VPWR final_adder.U$$469/X sky130_fd_sc_hd__a21o_1
XU$$308 U$$34/A1 U$$340/A2 U$$36/A1 U$$340/B2 VGND VGND VPWR VPWR U$$309/A sky130_fd_sc_hd__a22o_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$319 U$$319/A U$$353/B VGND VGND VPWR VPWR U$$319/X sky130_fd_sc_hd__xor2_1
XFILLER_38_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_112_1 U$$3689/X U$$3822/X U$$3955/X VGND VGND VPWR VPWR dadda_fa_4_113_1/CIN
+ dadda_fa_4_112_2/B sky130_fd_sc_hd__fa_1
XFILLER_153_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_105_0 U$$3675/X U$$3808/X U$$3941/X VGND VGND VPWR VPWR dadda_fa_4_106_0/B
+ dadda_fa_4_105_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_53_3 dadda_fa_3_53_3/A dadda_fa_3_53_3/B dadda_fa_3_53_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_1/B dadda_fa_4_53_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_69_3 U$$1608/X U$$1741/X U$$1874/X VGND VGND VPWR VPWR dadda_fa_1_70_7/A
+ dadda_fa_1_69_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_87_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_46_2 dadda_fa_3_46_2/A dadda_fa_3_46_2/B dadda_fa_3_46_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_1/A dadda_fa_4_46_2/B sky130_fd_sc_hd__fa_1
XFILLER_57_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$981 final_adder.U$$210/A final_adder.U$$823/X final_adder.U$$981/B1
+ VGND VGND VPWR VPWR final_adder.U$$981/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_3_39_1 dadda_fa_3_39_1/A dadda_fa_3_39_1/B dadda_fa_3_39_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_0/CIN dadda_fa_4_39_2/A sky130_fd_sc_hd__fa_1
XU$$820 U$$820/A U$$820/B VGND VGND VPWR VPWR U$$820/X sky130_fd_sc_hd__xor2_1
XU$$831 U$$831/A U$$875/B VGND VGND VPWR VPWR U$$831/X sky130_fd_sc_hd__xor2_1
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$842 U$$20/A1 U$$876/A2 U$$22/A1 U$$876/B2 VGND VGND VPWR VPWR U$$843/A sky130_fd_sc_hd__a22o_1
XU$$853 U$$853/A U$$907/B VGND VGND VPWR VPWR U$$853/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_16_0 dadda_fa_6_16_0/A dadda_fa_6_16_0/B dadda_fa_6_16_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_17_0/B dadda_fa_7_16_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1003 U$$44/A1 U$$979/A2 U$$46/A1 U$$979/B2 VGND VGND VPWR VPWR U$$1004/A sky130_fd_sc_hd__a22o_1
XU$$864 U$$864/A1 U$$898/A2 U$$864/B1 U$$898/B2 VGND VGND VPWR VPWR U$$865/A sky130_fd_sc_hd__a22o_1
XU$$1014 U$$1014/A U$$982/B VGND VGND VPWR VPWR U$$1014/X sky130_fd_sc_hd__xor2_1
XU$$875 U$$875/A U$$875/B VGND VGND VPWR VPWR U$$875/X sky130_fd_sc_hd__xor2_1
XU$$886 U$$64/A1 U$$902/A2 U$$66/A1 U$$902/B2 VGND VGND VPWR VPWR U$$887/A sky130_fd_sc_hd__a22o_1
XU$$1025 U$$64/B1 U$$997/A2 U$$66/B1 U$$997/B2 VGND VGND VPWR VPWR U$$1026/A sky130_fd_sc_hd__a22o_1
XU$$897 U$$897/A U$$925/B VGND VGND VPWR VPWR U$$897/X sky130_fd_sc_hd__xor2_1
XU$$1036 U$$1036/A U$$1062/B VGND VGND VPWR VPWR U$$1036/X sky130_fd_sc_hd__xor2_1
XU$$1047 U$$773/A1 U$$1093/A2 U$$773/B1 U$$1093/B2 VGND VGND VPWR VPWR U$$1048/A sky130_fd_sc_hd__a22o_1
XU$$1058 U$$1058/A U$$1062/B VGND VGND VPWR VPWR U$$1058/X sky130_fd_sc_hd__xor2_1
XU$$1069 U$$932/A1 U$$963/X U$$934/A1 U$$964/X VGND VGND VPWR VPWR U$$1070/A sky130_fd_sc_hd__a22o_1
XFILLER_32_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4491_1893 VGND VGND VPWR VPWR U$$4491_1893/HI U$$4491/B sky130_fd_sc_hd__conb_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1170 U$$4424/A1 VGND VGND VPWR VPWR U$$3189/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1181 U$$4011/A1 VGND VGND VPWR VPWR U$$447/B1 sky130_fd_sc_hd__buf_4
XFILLER_66_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1192 input70/X VGND VGND VPWR VPWR U$$4283/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_41_1 U$$1951/X U$$2084/X U$$2217/X VGND VGND VPWR VPWR dadda_fa_3_42_0/CIN
+ dadda_fa_3_41_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_82_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_34_0 U$$341/X U$$474/X U$$607/X VGND VGND VPWR VPWR dadda_fa_3_35_0/B
+ dadda_fa_3_34_2/B sky130_fd_sc_hd__fa_1
XFILLER_35_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2260 U$$68/A1 U$$2272/A2 U$$70/A1 U$$2272/B2 VGND VGND VPWR VPWR U$$2261/A sky130_fd_sc_hd__a22o_1
XFILLER_35_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2271 U$$2271/A U$$2273/B VGND VGND VPWR VPWR U$$2271/X sky130_fd_sc_hd__xor2_1
XU$$2282 U$$773/B1 U$$2282/A2 U$$640/A1 U$$2282/B2 VGND VGND VPWR VPWR U$$2283/A sky130_fd_sc_hd__a22o_1
XFILLER_34_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2293 U$$2293/A U$$2329/A VGND VGND VPWR VPWR U$$2293/X sky130_fd_sc_hd__xor2_1
XU$$1570 U$$1570/A U$$1570/B VGND VGND VPWR VPWR U$$1570/X sky130_fd_sc_hd__xor2_1
XU$$1581 U$$2814/A1 U$$1587/A2 U$$76/A1 U$$1587/B2 VGND VGND VPWR VPWR U$$1582/A sky130_fd_sc_hd__a22o_1
XU$$1592 U$$1592/A U$$1594/B VGND VGND VPWR VPWR U$$1592/X sky130_fd_sc_hd__xor2_1
XFILLER_31_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_86_3 U$$2706/X U$$2839/X U$$2972/X VGND VGND VPWR VPWR dadda_fa_2_87_3/CIN
+ dadda_fa_2_86_5/B sky130_fd_sc_hd__fa_1
XFILLER_103_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_63_2 dadda_fa_4_63_2/A dadda_fa_4_63_2/B dadda_fa_4_63_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_64_0/CIN dadda_fa_5_63_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_79_2 U$$1894/X U$$2027/X U$$2160/X VGND VGND VPWR VPWR dadda_fa_2_80_1/A
+ dadda_fa_2_79_4/A sky130_fd_sc_hd__fa_1
XFILLER_76_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_56_1 dadda_fa_4_56_1/A dadda_fa_4_56_1/B dadda_fa_4_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_57_0/B dadda_fa_5_56_1/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$200 final_adder.U$$200/A final_adder.U$$200/B VGND VGND VPWR VPWR
+ final_adder.U$$328/B sky130_fd_sc_hd__and2_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$211 final_adder.U$$210/B final_adder.U$$981/B1 final_adder.U$$211/B1
+ VGND VGND VPWR VPWR final_adder.U$$211/X sky130_fd_sc_hd__a21o_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_33_0 dadda_fa_7_33_0/A dadda_fa_7_33_0/B dadda_fa_7_33_0/CIN VGND VGND
+ VPWR VPWR _330_/D _201_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$222 final_adder.U$$222/A final_adder.U$$222/B VGND VGND VPWR VPWR
+ final_adder.U$$350/B sky130_fd_sc_hd__and2_1
Xdadda_fa_4_49_0 dadda_fa_4_49_0/A dadda_fa_4_49_0/B dadda_fa_4_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_50_0/A dadda_fa_5_49_1/A sky130_fd_sc_hd__fa_1
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$233 final_adder.U$$232/B final_adder.U$$233/A2 final_adder.U$$233/B1
+ VGND VGND VPWR VPWR final_adder.U$$233/X sky130_fd_sc_hd__a21o_1
XFILLER_58_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$244 final_adder.U$$244/A final_adder.U$$244/B VGND VGND VPWR VPWR
+ final_adder.U$$372/B sky130_fd_sc_hd__and2_1
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$255 final_adder.U$$1/SUM final_adder.U$$255/A2 final_adder.U$$255/B1
+ VGND VGND VPWR VPWR final_adder.U$$255/X sky130_fd_sc_hd__a21o_2
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$266 final_adder.U$$268/B final_adder.U$$266/B VGND VGND VPWR VPWR
+ final_adder.U$$392/B sky130_fd_sc_hd__and2_1
XU$$105 U$$105/A U$$127/B VGND VGND VPWR VPWR U$$105/X sky130_fd_sc_hd__xor2_1
XFILLER_85_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$277 final_adder.U$$276/B final_adder.U$$151/X final_adder.U$$149/X
+ VGND VGND VPWR VPWR final_adder.U$$277/X sky130_fd_sc_hd__a21o_1
XFILLER_73_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$116 U$$253/A1 U$$120/A2 U$$253/B1 U$$120/B2 VGND VGND VPWR VPWR U$$117/A sky130_fd_sc_hd__a22o_1
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$288 final_adder.U$$290/B final_adder.U$$288/B VGND VGND VPWR VPWR
+ final_adder.U$$414/B sky130_fd_sc_hd__and2_1
XU$$127 U$$127/A U$$127/B VGND VGND VPWR VPWR U$$127/X sky130_fd_sc_hd__xor2_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$299 final_adder.U$$298/B final_adder.U$$173/X final_adder.U$$171/X
+ VGND VGND VPWR VPWR final_adder.U$$299/X sky130_fd_sc_hd__a21o_1
XU$$138 U$$138/A VGND VGND VPWR VPWR U$$140/B sky130_fd_sc_hd__inv_1
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$149 U$$12/A1 U$$179/A2 U$$14/A1 U$$179/B2 VGND VGND VPWR VPWR U$$150/A sky130_fd_sc_hd__a22o_1
XFILLER_26_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_391_ _391_/CLK _391_/D VGND VGND VPWR VPWR _391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_clk _370_/CLK VGND VGND VPWR VPWR _421_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_74_1 U$$1086/X U$$1219/X U$$1352/X VGND VGND VPWR VPWR dadda_fa_1_75_8/A
+ dadda_fa_1_74_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput240 c[85] VGND VGND VPWR VPWR input240/X sky130_fd_sc_hd__dlymetal6s2s_1
Xdadda_fa_3_51_0 dadda_fa_3_51_0/A dadda_fa_3_51_0/B dadda_fa_3_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_0/B dadda_fa_4_51_1/CIN sky130_fd_sc_hd__fa_1
Xinput251 c[95] VGND VGND VPWR VPWR input251/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_0_67_0 U$$136/Y U$$273/Y U$$407/X VGND VGND VPWR VPWR dadda_fa_1_68_5/B
+ dadda_fa_1_67_7/B sky130_fd_sc_hd__fa_1
XFILLER_75_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$650 U$$650/A1 U$$682/A2 U$$650/B1 U$$682/B2 VGND VGND VPWR VPWR U$$651/A sky130_fd_sc_hd__a22o_1
XU$$661 U$$661/A U$$669/B VGND VGND VPWR VPWR U$$661/X sky130_fd_sc_hd__xor2_1
XU$$672 U$$672/A1 U$$676/A2 U$$672/B1 U$$676/B2 VGND VGND VPWR VPWR U$$673/A sky130_fd_sc_hd__a22o_1
XFILLER_90_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$683 U$$683/A U$$684/A VGND VGND VPWR VPWR U$$683/X sky130_fd_sc_hd__xor2_1
XU$$694 U$$694/A U$$744/B VGND VGND VPWR VPWR U$$694/X sky130_fd_sc_hd__xor2_1
XFILLER_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_11_clk _370_/CLK VGND VGND VPWR VPWR _247_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_118_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_96_2 U$$3258/X U$$3391/X U$$3524/X VGND VGND VPWR VPWR dadda_fa_3_97_1/A
+ dadda_fa_3_96_3/A sky130_fd_sc_hd__fa_1
XFILLER_173_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_73_1 dadda_fa_5_73_1/A dadda_fa_5_73_1/B dadda_fa_5_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_74_0/B dadda_fa_7_73_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_89_1 U$$3776/X U$$3909/X U$$4042/X VGND VGND VPWR VPWR dadda_fa_3_90_0/CIN
+ dadda_fa_3_89_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_98_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_66_0 dadda_fa_5_66_0/A dadda_fa_5_66_0/B dadda_fa_5_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_67_0/A dadda_fa_6_66_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_63_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout407 U$$689/X VGND VGND VPWR VPWR U$$819/A2 sky130_fd_sc_hd__buf_4
XFILLER_99_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout418 U$$4309/A2 VGND VGND VPWR VPWR U$$4381/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_98_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout429 U$$545/A2 VGND VGND VPWR VPWR U$$447/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_65_8 dadda_fa_1_65_8/A dadda_fa_1_65_8/B dadda_fa_1_65_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_66_3/A dadda_fa_3_65_0/A sky130_fd_sc_hd__fa_2
XFILLER_79_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_58_7 dadda_fa_1_58_7/A dadda_fa_1_58_7/B dadda_fa_1_58_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_59_2/CIN dadda_fa_2_58_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_54_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_858 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_5_0 U$$283/X input212/X dadda_fa_6_5_0/CIN VGND VGND VPWR VPWR dadda_fa_7_6_0/B
+ dadda_fa_7_5_0/CIN sky130_fd_sc_hd__fa_1
XU$$2090 U$$2090/A U$$2096/B VGND VGND VPWR VPWR U$$2090/X sky130_fd_sc_hd__xor2_1
XFILLER_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_91_1 U$$2317/X U$$2450/X U$$2583/X VGND VGND VPWR VPWR dadda_fa_2_92_4/CIN
+ dadda_fa_2_91_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_151_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_84_0 dadda_fa_1_84_0/A U$$1505/X U$$1638/X VGND VGND VPWR VPWR dadda_fa_2_85_2/A
+ dadda_fa_2_84_4/A sky130_fd_sc_hd__fa_1
XFILLER_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout930 fanout938/X VGND VGND VPWR VPWR U$$88/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_89_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout941 U$$4259/B1 VGND VGND VPWR VPWR U$$2480/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout952 fanout957/X VGND VGND VPWR VPWR U$$3509/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_77_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout963 fanout966/X VGND VGND VPWR VPWR U$$3920/A1 sky130_fd_sc_hd__buf_2
XFILLER_93_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4409 U$$4409/A U$$4409/B VGND VGND VPWR VPWR U$$4409/X sky130_fd_sc_hd__xor2_1
XFILLER_161_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout974 fanout975/X VGND VGND VPWR VPWR U$$4466/A1 sky130_fd_sc_hd__buf_4
Xfanout985 fanout993/X VGND VGND VPWR VPWR U$$900/A1 sky130_fd_sc_hd__buf_4
Xfanout996 U$$3775/A1 VGND VGND VPWR VPWR U$$3636/B1 sky130_fd_sc_hd__buf_4
XFILLER_58_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3708 U$$3708/A U$$3790/B VGND VGND VPWR VPWR U$$3708/X sky130_fd_sc_hd__xor2_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3719 U$$4265/B1 U$$3757/A2 U$$4132/A1 U$$3757/B2 VGND VGND VPWR VPWR U$$3720/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_374_ _375_/CLK _374_/D VGND VGND VPWR VPWR _374_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4403_1849 VGND VGND VPWR VPWR U$$4403_1849/HI U$$4403/B sky130_fd_sc_hd__conb_1
XFILLER_174_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_83_0 dadda_fa_6_83_0/A dadda_fa_6_83_0/B dadda_fa_6_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_84_0/B dadda_fa_7_83_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_154_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_99_0 U$$4461/X input255/X dadda_fa_3_99_0/CIN VGND VGND VPWR VPWR dadda_fa_4_100_0/B
+ dadda_fa_4_99_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_clk _201_/CLK VGND VGND VPWR VPWR _349_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$480 U$$480/A U$$480/B VGND VGND VPWR VPWR U$$480/X sky130_fd_sc_hd__xor2_1
XU$$491 U$$900/B1 U$$497/A2 U$$765/B1 U$$497/B2 VGND VGND VPWR VPWR U$$492/A sky130_fd_sc_hd__a22o_1
XFILLER_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_70_6 dadda_fa_1_70_6/A dadda_fa_1_70_6/B dadda_fa_1_70_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_71_2/B dadda_fa_2_70_5/B sky130_fd_sc_hd__fa_1
XFILLER_86_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_63_5 input216/X dadda_fa_1_63_5/B dadda_fa_1_63_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_64_2/A dadda_fa_2_63_5/A sky130_fd_sc_hd__fa_1
XFILLER_75_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_56_4 U$$2779/X U$$2912/X U$$3045/X VGND VGND VPWR VPWR dadda_fa_2_57_1/CIN
+ dadda_fa_2_56_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_49_3 U$$1302/X U$$1435/X U$$1568/X VGND VGND VPWR VPWR dadda_fa_2_50_1/CIN
+ dadda_fa_2_49_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_82_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_26_2 dadda_fa_4_26_2/A dadda_fa_4_26_2/B dadda_fa_4_26_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_27_0/CIN dadda_fa_5_26_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_19_1 dadda_fa_4_19_1/A dadda_fa_4_19_1/B dadda_fa_4_19_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_20_0/B dadda_fa_5_19_1/B sky130_fd_sc_hd__fa_1
XFILLER_23_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_922 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1703 fanout1708/X VGND VGND VPWR VPWR U$$654/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout1714 fanout1718/X VGND VGND VPWR VPWR U$$650/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1725 U$$4486/A1 VGND VGND VPWR VPWR U$$4484/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1736 U$$370/B1 VGND VGND VPWR VPWR U$$2973/B1 sky130_fd_sc_hd__buf_4
XFILLER_131_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1747 input103/X VGND VGND VPWR VPWR U$$505/B1 sky130_fd_sc_hd__buf_6
XFILLER_133_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout760 U$$3293/X VGND VGND VPWR VPWR U$$3306/B2 sky130_fd_sc_hd__buf_4
XU$$4206 U$$4480/A1 U$$4226/A2 U$$4482/A1 U$$4226/B2 VGND VGND VPWR VPWR U$$4207/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1758 U$$3382/A1 VGND VGND VPWR VPWR U$$4478/A1 sky130_fd_sc_hd__buf_4
Xfanout771 U$$3112/B2 VGND VGND VPWR VPWR U$$3072/B2 sky130_fd_sc_hd__buf_4
XU$$4217 U$$4217/A U$$4231/B VGND VGND VPWR VPWR U$$4217/X sky130_fd_sc_hd__xor2_1
Xfanout1769 U$$914/A1 VGND VGND VPWR VPWR U$$3515/B1 sky130_fd_sc_hd__buf_4
Xfanout782 U$$2882/X VGND VGND VPWR VPWR U$$2977/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4228 U$$4365/A1 U$$4236/A2 U$$4365/B1 U$$4236/B2 VGND VGND VPWR VPWR U$$4229/A
+ sky130_fd_sc_hd__a22o_1
XU$$4239 U$$4239/A U$$4241/B VGND VGND VPWR VPWR U$$4239/X sky130_fd_sc_hd__xor2_1
Xfanout793 U$$338/B2 VGND VGND VPWR VPWR U$$346/B2 sky130_fd_sc_hd__clkbuf_2
XU$$3505 U$$3642/A1 U$$3505/A2 U$$3642/B1 U$$3505/B2 VGND VGND VPWR VPWR U$$3506/A
+ sky130_fd_sc_hd__a22o_1
XU$$3516 U$$3516/A U$$3558/B VGND VGND VPWR VPWR U$$3516/X sky130_fd_sc_hd__xor2_1
XU$$3527 U$$4349/A1 U$$3549/A2 U$$4349/B1 U$$3549/B2 VGND VGND VPWR VPWR U$$3528/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3538 U$$3538/A U$$3548/B VGND VGND VPWR VPWR U$$3538/X sky130_fd_sc_hd__xor2_1
XU$$2804 U$$3763/A1 U$$2804/A2 U$$3628/A1 U$$2804/B2 VGND VGND VPWR VPWR U$$2805/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3549 U$$3684/B1 U$$3549/A2 U$$3551/A1 U$$3549/B2 VGND VGND VPWR VPWR U$$3550/A
+ sky130_fd_sc_hd__a22o_1
XU$$2815 U$$2815/A U$$2873/B VGND VGND VPWR VPWR U$$2815/X sky130_fd_sc_hd__xor2_1
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2826 U$$3372/B1 U$$2840/A2 U$$3239/A1 U$$2840/B2 VGND VGND VPWR VPWR U$$2827/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2837 U$$2837/A U$$2841/B VGND VGND VPWR VPWR U$$2837/X sky130_fd_sc_hd__xor2_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2848 U$$4353/B1 U$$2874/A2 U$$4220/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2849/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_21_1 U$$448/X U$$581/X U$$714/X VGND VGND VPWR VPWR dadda_fa_4_22_0/CIN
+ dadda_fa_4_21_2/A sky130_fd_sc_hd__fa_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2859 U$$2859/A U$$2871/B VGND VGND VPWR VPWR U$$2859/X sky130_fd_sc_hd__xor2_1
XFILLER_61_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_357_ _358_/CLK _357_/D VGND VGND VPWR VPWR _357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_288_ _421_/CLK _288_/D VGND VGND VPWR VPWR _288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_80_5 dadda_fa_2_80_5/A dadda_fa_2_80_5/B dadda_fa_2_80_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_2/A dadda_fa_4_80_0/A sky130_fd_sc_hd__fa_2
XFILLER_114_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_73_4 dadda_fa_2_73_4/A dadda_fa_2_73_4/B dadda_fa_2_73_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_1/CIN dadda_fa_3_73_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_66_3 dadda_fa_2_66_3/A dadda_fa_2_66_3/B dadda_fa_2_66_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_1/B dadda_fa_3_66_3/B sky130_fd_sc_hd__fa_1
XFILLER_57_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_59_2 dadda_fa_2_59_2/A dadda_fa_2_59_2/B dadda_fa_2_59_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_1/A dadda_fa_3_59_3/A sky130_fd_sc_hd__fa_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput4 a[12] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_5_36_1 dadda_fa_5_36_1/A dadda_fa_5_36_1/B dadda_fa_5_36_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_37_0/B dadda_fa_7_36_0/A sky130_fd_sc_hd__fa_1
XFILLER_65_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_29_0 dadda_fa_5_29_0/A dadda_fa_5_29_0/B dadda_fa_5_29_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_30_0/A dadda_fa_6_29_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_25_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1__f_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _201_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_956 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4425_1860 VGND VGND VPWR VPWR U$$4425_1860/HI U$$4425/B sky130_fd_sc_hd__conb_1
XFILLER_20_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_110_1 dadda_fa_5_110_1/A dadda_fa_5_110_1/B dadda_fa_5_110_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_111_0/B dadda_fa_7_110_0/A sky130_fd_sc_hd__fa_1
XFILLER_119_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$2 _298_/Q _170_/Q VGND VGND VPWR VPWR final_adder.U$$253/A2 final_adder.U$$252/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_5_103_0 dadda_fa_5_103_0/A dadda_fa_5_103_0/B dadda_fa_5_103_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_104_0/A dadda_fa_6_103_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput330 output330/A VGND VGND VPWR VPWR o[50] sky130_fd_sc_hd__buf_2
Xoutput341 output341/A VGND VGND VPWR VPWR o[60] sky130_fd_sc_hd__buf_2
XFILLER_160_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput352 output352/A VGND VGND VPWR VPWR o[70] sky130_fd_sc_hd__buf_2
Xoutput363 output363/A VGND VGND VPWR VPWR o[80] sky130_fd_sc_hd__buf_2
Xoutput374 output374/A VGND VGND VPWR VPWR o[90] sky130_fd_sc_hd__buf_2
XFILLER_99_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3148_1815 VGND VGND VPWR VPWR U$$3148_1815/HI U$$3148/B1 sky130_fd_sc_hd__conb_1
XFILLER_99_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_61_2 U$$2789/X U$$2922/X U$$3055/X VGND VGND VPWR VPWR dadda_fa_2_62_1/A
+ dadda_fa_2_61_4/A sky130_fd_sc_hd__fa_1
XFILLER_101_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_1 U$$1179/X U$$1312/X U$$1445/X VGND VGND VPWR VPWR dadda_fa_2_55_0/CIN
+ dadda_fa_2_54_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_19_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_31_0 dadda_fa_4_31_0/A dadda_fa_4_31_0/B dadda_fa_4_31_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_32_0/A dadda_fa_5_31_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_47_0 U$$101/X U$$234/X U$$367/X VGND VGND VPWR VPWR dadda_fa_2_48_1/B
+ dadda_fa_2_47_4/A sky130_fd_sc_hd__fa_1
XFILLER_27_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_211_ _346_/CLK _211_/D VGND VGND VPWR VPWR _211_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_83_3 dadda_fa_3_83_3/A dadda_fa_3_83_3/B dadda_fa_3_83_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_1/B dadda_fa_4_83_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_76_2 dadda_fa_3_76_2/A dadda_fa_3_76_2/B dadda_fa_3_76_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_1/A dadda_fa_4_76_2/B sky130_fd_sc_hd__fa_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1500 U$$1455/B VGND VGND VPWR VPWR U$$1449/B sky130_fd_sc_hd__buf_8
Xdadda_fa_3_69_1 dadda_fa_3_69_1/A dadda_fa_3_69_1/B dadda_fa_3_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_0/CIN dadda_fa_4_69_2/A sky130_fd_sc_hd__fa_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1511 U$$3314/A1 VGND VGND VPWR VPWR U$$26/A1 sky130_fd_sc_hd__buf_4
Xfanout1522 input127/X VGND VGND VPWR VPWR U$$4408/A1 sky130_fd_sc_hd__buf_4
Xfanout1533 U$$4404/A1 VGND VGND VPWR VPWR U$$4265/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_6_46_0 dadda_fa_6_46_0/A dadda_fa_6_46_0/B dadda_fa_6_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_47_0/B dadda_fa_7_46_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_116_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1544 U$$3559/A1 VGND VGND VPWR VPWR U$$3833/A1 sky130_fd_sc_hd__buf_2
XU$$4003 U$$987/B1 U$$4005/A2 input68/X U$$4005/B2 VGND VGND VPWR VPWR U$$4004/A sky130_fd_sc_hd__a22o_1
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1555 input123/X VGND VGND VPWR VPWR U$$954/A1 sky130_fd_sc_hd__buf_4
Xfanout1566 U$$4512/A1 VGND VGND VPWR VPWR U$$811/B1 sky130_fd_sc_hd__buf_2
XU$$4014 U$$4014/A U$$4058/B VGND VGND VPWR VPWR U$$4014/X sky130_fd_sc_hd__xor2_1
Xfanout1577 input120/X VGND VGND VPWR VPWR U$$4402/A1 sky130_fd_sc_hd__buf_4
XU$$4025 U$$4162/A1 U$$4025/A2 U$$4162/B1 U$$4025/B2 VGND VGND VPWR VPWR U$$4026/A
+ sky130_fd_sc_hd__a22o_1
XU$$4036 U$$4036/A U$$4040/B VGND VGND VPWR VPWR U$$4036/X sky130_fd_sc_hd__xor2_1
Xfanout590 U$$2052/A2 VGND VGND VPWR VPWR U$$2046/A2 sky130_fd_sc_hd__buf_4
Xfanout1588 U$$81/B VGND VGND VPWR VPWR U$$49/B sky130_fd_sc_hd__clkbuf_4
XU$$3302 U$$562/A1 U$$3306/A2 U$$562/B1 U$$3306/B2 VGND VGND VPWR VPWR U$$3303/A sky130_fd_sc_hd__a22o_1
Xfanout1599 U$$2729/A1 VGND VGND VPWR VPWR U$$3960/B1 sky130_fd_sc_hd__clkbuf_2
XU$$4047 U$$4458/A1 U$$4105/A2 U$$4049/A1 U$$4105/B2 VGND VGND VPWR VPWR U$$4048/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3313 U$$3313/A U$$3349/B VGND VGND VPWR VPWR U$$3313/X sky130_fd_sc_hd__xor2_1
XU$$4058 U$$4058/A U$$4058/B VGND VGND VPWR VPWR U$$4058/X sky130_fd_sc_hd__xor2_1
XU$$3324 U$$3870/B1 U$$3338/A2 U$$4420/B1 U$$3338/B2 VGND VGND VPWR VPWR U$$3325/A
+ sky130_fd_sc_hd__a22o_1
XU$$4069 U$$4480/A1 U$$4081/A2 U$$4482/A1 U$$4081/B2 VGND VGND VPWR VPWR U$$4070/A
+ sky130_fd_sc_hd__a22o_1
XU$$3335 U$$3335/A U$$3335/B VGND VGND VPWR VPWR U$$3335/X sky130_fd_sc_hd__xor2_1
XU$$2601 U$$2601/A U$$2602/A VGND VGND VPWR VPWR U$$2601/X sky130_fd_sc_hd__xor2_1
XU$$3346 U$$3618/B1 U$$3390/A2 U$$4444/A1 U$$3390/B2 VGND VGND VPWR VPWR U$$3347/A
+ sky130_fd_sc_hd__a22o_1
XU$$2612 U$$2612/A U$$2678/B VGND VGND VPWR VPWR U$$2612/X sky130_fd_sc_hd__xor2_1
XU$$3357 U$$3357/A U$$3373/B VGND VGND VPWR VPWR U$$3357/X sky130_fd_sc_hd__xor2_1
XFILLER_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_105_2 dadda_fa_4_105_2/A dadda_fa_4_105_2/B dadda_fa_4_105_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_106_0/CIN dadda_fa_5_105_1/CIN sky130_fd_sc_hd__fa_1
XU$$2623 U$$2758/B1 U$$2665/A2 U$$2625/A1 U$$2665/B2 VGND VGND VPWR VPWR U$$2624/A
+ sky130_fd_sc_hd__a22o_1
XU$$3368 U$$3503/B1 U$$3372/A2 U$$3370/A1 U$$3372/B2 VGND VGND VPWR VPWR U$$3369/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3379 U$$3379/A U$$3425/A VGND VGND VPWR VPWR U$$3379/X sky130_fd_sc_hd__xor2_1
XU$$2634 U$$2634/A U$$2678/B VGND VGND VPWR VPWR U$$2634/X sky130_fd_sc_hd__xor2_1
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1900 U$$1900/A U$$1910/B VGND VGND VPWR VPWR U$$1900/X sky130_fd_sc_hd__xor2_1
XU$$2645 U$$2780/B1 U$$2681/A2 U$$44/A1 U$$2681/B2 VGND VGND VPWR VPWR U$$2646/A sky130_fd_sc_hd__a22o_1
XU$$1911 U$$4512/B1 U$$1911/A2 U$$4377/B1 U$$1911/B2 VGND VGND VPWR VPWR U$$1912/A
+ sky130_fd_sc_hd__a22o_1
XU$$2656 U$$2656/A U$$2662/B VGND VGND VPWR VPWR U$$2656/X sky130_fd_sc_hd__xor2_1
XU$$1922 U$$1920/Y input21/X U$$1918/A U$$1921/X U$$1918/Y VGND VGND VPWR VPWR U$$1922/X
+ sky130_fd_sc_hd__a32o_1
XU$$2667 U$$3763/A1 U$$2667/A2 U$$3628/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2668/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1933 U$$1933/A U$$1971/B VGND VGND VPWR VPWR U$$1933/X sky130_fd_sc_hd__xor2_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2678 U$$2678/A U$$2678/B VGND VGND VPWR VPWR U$$2678/X sky130_fd_sc_hd__xor2_1
XFILLER_62_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2689 U$$4470/A1 U$$2711/A2 U$$3650/A1 U$$2711/B2 VGND VGND VPWR VPWR U$$2690/A
+ sky130_fd_sc_hd__a22o_1
XU$$1944 U$$709/B1 U$$1986/A2 U$$576/A1 U$$1986/B2 VGND VGND VPWR VPWR U$$1945/A sky130_fd_sc_hd__a22o_1
XU$$1955 U$$1955/A U$$1963/B VGND VGND VPWR VPWR U$$1955/X sky130_fd_sc_hd__xor2_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1966 U$$2925/A1 U$$1986/A2 U$$735/A1 U$$1986/B2 VGND VGND VPWR VPWR U$$1967/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1977 U$$1977/A U$$1981/B VGND VGND VPWR VPWR U$$1977/X sky130_fd_sc_hd__xor2_1
XFILLER_30_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1988 U$$70/A1 U$$2006/A2 U$$70/B1 U$$2006/B2 VGND VGND VPWR VPWR U$$1989/A sky130_fd_sc_hd__a22o_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1999 U$$1999/A U$$2031/B VGND VGND VPWR VPWR U$$1999/X sky130_fd_sc_hd__xor2_1
X_409_ _416_/CLK _409_/D VGND VGND VPWR VPWR _409_/Q sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_7_119_0 dadda_fa_7_119_0/A dadda_fa_7_119_0/B dadda_fa_7_119_0/CIN VGND
+ VGND VPWR VPWR _416_/D _287_/D sky130_fd_sc_hd__fa_1
XFILLER_174_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4455_1875 VGND VGND VPWR VPWR U$$4455_1875/HI U$$4455/B sky130_fd_sc_hd__conb_1
XFILLER_170_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_71_1 dadda_fa_2_71_1/A dadda_fa_2_71_1/B dadda_fa_2_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_0/CIN dadda_fa_3_71_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_97_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_64_0 dadda_fa_2_64_0/A dadda_fa_2_64_0/B dadda_fa_2_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_0/B dadda_fa_3_64_2/B sky130_fd_sc_hd__fa_1
XFILLER_97_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$607 final_adder.U$$606/B final_adder.U$$491/X final_adder.U$$483/X
+ VGND VGND VPWR VPWR final_adder.U$$607/X sky130_fd_sc_hd__a21o_1
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$629 final_adder.U$$628/B final_adder.U$$525/X final_adder.U$$509/X
+ VGND VGND VPWR VPWR final_adder.U$$629/X sky130_fd_sc_hd__a21o_1
XFILLER_56_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$40 U$$40/A1 U$$74/A2 U$$40/B1 U$$74/B2 VGND VGND VPWR VPWR U$$41/A sky130_fd_sc_hd__a22o_1
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$51 U$$51/A U$$87/B VGND VGND VPWR VPWR U$$51/X sky130_fd_sc_hd__xor2_1
XU$$62 U$$62/A1 U$$96/A2 U$$64/A1 U$$96/B2 VGND VGND VPWR VPWR U$$63/A sky130_fd_sc_hd__a22o_1
XFILLER_25_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$73 U$$73/A U$$77/B VGND VGND VPWR VPWR U$$73/X sky130_fd_sc_hd__xor2_1
XFILLER_53_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$84 U$$84/A1 U$$86/A2 U$$86/A1 U$$86/B2 VGND VGND VPWR VPWR U$$85/A sky130_fd_sc_hd__a22o_1
XU$$3880 U$$4152/B1 U$$3924/A2 U$$4017/B1 U$$3924/B2 VGND VGND VPWR VPWR U$$3881/A
+ sky130_fd_sc_hd__a22o_1
XU$$3891 U$$3891/A U$$3907/B VGND VGND VPWR VPWR U$$3891/X sky130_fd_sc_hd__xor2_1
XFILLER_24_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$95 U$$95/A U$$97/B VGND VGND VPWR VPWR U$$95/X sky130_fd_sc_hd__xor2_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_93_2 dadda_fa_4_93_2/A dadda_fa_4_93_2/B dadda_fa_4_93_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_94_0/CIN dadda_fa_5_93_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_86_1 dadda_fa_4_86_1/A dadda_fa_4_86_1/B dadda_fa_4_86_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_87_0/B dadda_fa_5_86_1/B sky130_fd_sc_hd__fa_1
XFILLER_118_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_63_0 dadda_fa_7_63_0/A dadda_fa_7_63_0/B dadda_fa_7_63_0/CIN VGND VGND
+ VPWR VPWR _360_/D _231_/D sky130_fd_sc_hd__fa_1
XFILLER_106_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_79_0 dadda_fa_4_79_0/A dadda_fa_4_79_0/B dadda_fa_4_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_80_0/A dadda_fa_5_79_1/A sky130_fd_sc_hd__fa_1
XFILLER_133_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_80_0_1923 VGND VGND VPWR VPWR dadda_fa_1_80_0/A dadda_fa_1_80_0_1923/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1207 U$$1207/A U$$1231/B VGND VGND VPWR VPWR U$$1207/X sky130_fd_sc_hd__xor2_1
XU$$1218 U$$120/B1 U$$1218/A2 U$$946/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1219/A sky130_fd_sc_hd__a22o_1
XFILLER_16_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1229 U$$1229/A U$$1231/B VGND VGND VPWR VPWR U$$1229/X sky130_fd_sc_hd__xor2_1
XFILLER_70_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1001 final_adder.U$$230/A final_adder.U$$731/X final_adder.U$$231/A2
+ VGND VGND VPWR VPWR final_adder.U$$1049/B sky130_fd_sc_hd__a21o_1
XFILLER_157_858 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$1023 final_adder.U$$252/A final_adder.U$$255/X final_adder.U$$253/A2
+ VGND VGND VPWR VPWR final_adder.U$$1027/B sky130_fd_sc_hd__a21o_1
XFILLER_7_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1034 final_adder.U$$244/A final_adder.U$$625/X VGND VGND VPWR VPWR
+ output268/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1045 final_adder.U$$234/B final_adder.U$$1045/B VGND VGND VPWR VPWR
+ output298/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1056 final_adder.U$$222/A final_adder.U$$723/X VGND VGND VPWR VPWR
+ output310/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1067 final_adder.U$$212/B final_adder.U$$983/X VGND VGND VPWR VPWR
+ output322/A sky130_fd_sc_hd__xor2_1
XFILLER_7_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1078 final_adder.U$$200/A final_adder.U$$813/X VGND VGND VPWR VPWR
+ output334/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1089 final_adder.U$$190/B final_adder.U$$961/X VGND VGND VPWR VPWR
+ output346/A sky130_fd_sc_hd__xor2_1
XFILLER_152_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_81_0 dadda_fa_3_81_0/A dadda_fa_3_81_0/B dadda_fa_3_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_0/B dadda_fa_4_81_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1330 U$$3607/B VGND VGND VPWR VPWR U$$3699/A sky130_fd_sc_hd__buf_4
XFILLER_87_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1341 U$$3524/B VGND VGND VPWR VPWR U$$3482/B sky130_fd_sc_hd__buf_6
XFILLER_78_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1352 U$$3424/A VGND VGND VPWR VPWR U$$3411/B sky130_fd_sc_hd__buf_2
Xfanout1363 fanout1364/X VGND VGND VPWR VPWR U$$3287/A sky130_fd_sc_hd__buf_4
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1374 U$$2938/B VGND VGND VPWR VPWR U$$2926/B sky130_fd_sc_hd__buf_4
XFILLER_94_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1385 fanout1391/X VGND VGND VPWR VPWR U$$2841/B sky130_fd_sc_hd__buf_6
Xfanout1396 input34/X VGND VGND VPWR VPWR U$$260/B sky130_fd_sc_hd__buf_6
XU$$3110 U$$3110/A1 U$$3112/A2 U$$3112/A1 U$$3112/B2 VGND VGND VPWR VPWR U$$3111/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_43_5 dadda_fa_2_43_5/A dadda_fa_2_43_5/B dadda_fa_2_43_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_44_2/A dadda_fa_4_43_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_4_110_0 input141/X dadda_fa_4_110_0/B dadda_fa_4_110_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_5_111_0/A dadda_fa_5_110_1/A sky130_fd_sc_hd__fa_1
XU$$3121 U$$3121/A U$$3150/A VGND VGND VPWR VPWR U$$3121/X sky130_fd_sc_hd__xor2_1
XU$$3132 U$$3817/A1 U$$3144/A2 U$$3817/B1 U$$3144/B2 VGND VGND VPWR VPWR U$$3133/A
+ sky130_fd_sc_hd__a22o_1
XU$$3143 U$$3143/A U$$3147/B VGND VGND VPWR VPWR U$$3143/X sky130_fd_sc_hd__xor2_1
XFILLER_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3154 U$$3288/A U$$3154/B VGND VGND VPWR VPWR U$$3154/X sky130_fd_sc_hd__and2_1
XFILLER_62_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3165 U$$973/A1 U$$3255/A2 U$$973/B1 U$$3255/B2 VGND VGND VPWR VPWR U$$3166/A sky130_fd_sc_hd__a22o_1
XU$$2420 U$$2420/A U$$2456/B VGND VGND VPWR VPWR U$$2420/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_36_4 U$$2340/X U$$2473/X U$$2549/B VGND VGND VPWR VPWR dadda_fa_3_37_1/CIN
+ dadda_fa_3_36_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2431 U$$2840/B1 U$$2443/A2 U$$2707/A1 U$$2443/B2 VGND VGND VPWR VPWR U$$2432/A
+ sky130_fd_sc_hd__a22o_1
XU$$3176 U$$3176/A U$$3210/B VGND VGND VPWR VPWR U$$3176/X sky130_fd_sc_hd__xor2_1
XU$$2442 U$$2442/A U$$2466/A VGND VGND VPWR VPWR U$$2442/X sky130_fd_sc_hd__xor2_1
XU$$3187 U$$3322/B1 U$$3199/A2 U$$3189/A1 U$$3199/B2 VGND VGND VPWR VPWR U$$3188/A
+ sky130_fd_sc_hd__a22o_1
XU$$3198 U$$3198/A U$$3208/B VGND VGND VPWR VPWR U$$3198/X sky130_fd_sc_hd__xor2_1
XU$$2453 U$$4234/A1 U$$2459/A2 U$$4234/B1 U$$2459/B2 VGND VGND VPWR VPWR U$$2454/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2464 U$$2464/A U$$2465/A VGND VGND VPWR VPWR U$$2464/X sky130_fd_sc_hd__xor2_1
XU$$1730 U$$3372/B1 U$$1774/A2 U$$3239/A1 U$$1774/B2 VGND VGND VPWR VPWR U$$1731/A
+ sky130_fd_sc_hd__a22o_1
XU$$2475 U$$2475/A U$$2545/B VGND VGND VPWR VPWR U$$2475/X sky130_fd_sc_hd__xor2_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2486 U$$2758/B1 U$$2532/A2 U$$2625/A1 U$$2532/B2 VGND VGND VPWR VPWR U$$2487/A
+ sky130_fd_sc_hd__a22o_1
XU$$1741 U$$1741/A U$$1741/B VGND VGND VPWR VPWR U$$1741/X sky130_fd_sc_hd__xor2_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1752 U$$4353/B1 U$$1758/A2 U$$4220/A1 U$$1758/B2 VGND VGND VPWR VPWR U$$1753/A
+ sky130_fd_sc_hd__a22o_1
XU$$2497 U$$2497/A U$$2541/B VGND VGND VPWR VPWR U$$2497/X sky130_fd_sc_hd__xor2_1
XFILLER_61_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1763 U$$1763/A U$$1777/B VGND VGND VPWR VPWR U$$1763/X sky130_fd_sc_hd__xor2_1
XU$$1774 U$$4512/B1 U$$1774/A2 U$$4377/B1 U$$1774/B2 VGND VGND VPWR VPWR U$$1775/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1785 U$$1783/Y input19/X U$$1741/B U$$1784/X U$$1781/Y VGND VGND VPWR VPWR U$$1785/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_148_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1796 U$$1796/A U$$1832/B VGND VGND VPWR VPWR U$$1796/X sky130_fd_sc_hd__xor2_1
XFILLER_148_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_96_0 dadda_fa_5_96_0/A dadda_fa_5_96_0/B dadda_fa_5_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_97_0/A dadda_fa_6_96_0/CIN sky130_fd_sc_hd__fa_1
Xinput40 a[45] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__buf_4
XFILLER_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput51 a[55] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_1
Xinput62 a[7] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_2
Xinput73 b[17] VGND VGND VPWR VPWR input73/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput84 b[27] VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__buf_6
Xinput95 b[37] VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$404 final_adder.U$$408/B final_adder.U$$404/B VGND VGND VPWR VPWR
+ final_adder.U$$528/B sky130_fd_sc_hd__and2_1
XFILLER_29_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$415 final_adder.U$$414/B final_adder.U$$293/X final_adder.U$$289/X
+ VGND VGND VPWR VPWR final_adder.U$$415/X sky130_fd_sc_hd__a21o_1
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$426 final_adder.U$$430/B final_adder.U$$426/B VGND VGND VPWR VPWR
+ final_adder.U$$550/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$437 final_adder.U$$436/B final_adder.U$$315/X final_adder.U$$311/X
+ VGND VGND VPWR VPWR final_adder.U$$437/X sky130_fd_sc_hd__a21o_1
XFILLER_111_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$448 final_adder.U$$452/B final_adder.U$$448/B VGND VGND VPWR VPWR
+ final_adder.U$$572/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$459 final_adder.U$$458/B final_adder.U$$337/X final_adder.U$$333/X
+ VGND VGND VPWR VPWR final_adder.U$$459/X sky130_fd_sc_hd__a21o_1
XFILLER_26_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$309 U$$309/A U$$339/B VGND VGND VPWR VPWR U$$309/X sky130_fd_sc_hd__xor2_1
XFILLER_84_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_105_1 U$$4074/X U$$4207/X U$$4340/X VGND VGND VPWR VPWR dadda_fa_4_106_0/CIN
+ dadda_fa_4_105_2/A sky130_fd_sc_hd__fa_1
XFILLER_164_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_126_0 U$$4515/X input158/X dadda_fa_6_126_0/CIN VGND VGND VPWR VPWR dadda_fa_7_127_0/B
+ dadda_fa_7_126_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_69_4 U$$2007/X U$$2140/X U$$2273/X VGND VGND VPWR VPWR dadda_fa_1_70_7/B
+ dadda_fa_2_69_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_46_3 dadda_fa_3_46_3/A dadda_fa_3_46_3/B dadda_fa_3_46_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_1/B dadda_fa_4_46_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_169_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$971 final_adder.U$$200/A final_adder.U$$813/X final_adder.U$$971/B1
+ VGND VGND VPWR VPWR final_adder.U$$971/X sky130_fd_sc_hd__a21o_1
XFILLER_63_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$810 U$$810/A U$$822/A VGND VGND VPWR VPWR U$$810/X sky130_fd_sc_hd__xor2_1
XFILLER_90_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_39_2 dadda_fa_3_39_2/A dadda_fa_3_39_2/B dadda_fa_3_39_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_1/A dadda_fa_4_39_2/B sky130_fd_sc_hd__fa_1
XU$$821 U$$821/A VGND VGND VPWR VPWR U$$821/Y sky130_fd_sc_hd__inv_1
XFILLER_17_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$993 final_adder.U$$222/A final_adder.U$$723/X final_adder.U$$993/B1
+ VGND VGND VPWR VPWR final_adder.U$$993/X sky130_fd_sc_hd__a21o_1
XFILLER_56_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$832 U$$10/A1 U$$876/A2 U$$12/A1 U$$876/B2 VGND VGND VPWR VPWR U$$833/A sky130_fd_sc_hd__a22o_1
XU$$843 U$$843/A U$$875/B VGND VGND VPWR VPWR U$$843/X sky130_fd_sc_hd__xor2_1
XU$$854 U$$854/A1 U$$902/A2 U$$854/B1 U$$902/B2 VGND VGND VPWR VPWR U$$855/A sky130_fd_sc_hd__a22o_1
XU$$865 U$$865/A U$$895/B VGND VGND VPWR VPWR U$$865/X sky130_fd_sc_hd__xor2_1
XFILLER_90_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1004 U$$1004/A U$$980/B VGND VGND VPWR VPWR U$$1004/X sky130_fd_sc_hd__xor2_1
XU$$1015 U$$741/A1 U$$981/A2 U$$880/A1 U$$981/B2 VGND VGND VPWR VPWR U$$1016/A sky130_fd_sc_hd__a22o_1
XU$$876 U$$876/A1 U$$876/A2 U$$878/A1 U$$876/B2 VGND VGND VPWR VPWR U$$877/A sky130_fd_sc_hd__a22o_1
XU$$1026 U$$1026/A U$$998/B VGND VGND VPWR VPWR U$$1026/X sky130_fd_sc_hd__xor2_1
XU$$887 U$$887/A U$$925/B VGND VGND VPWR VPWR U$$887/X sky130_fd_sc_hd__xor2_1
XFILLER_43_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$898 U$$898/A1 U$$898/A2 U$$900/A1 U$$898/B2 VGND VGND VPWR VPWR U$$899/A sky130_fd_sc_hd__a22o_1
XU$$1037 U$$215/A1 U$$981/A2 U$$215/B1 U$$981/B2 VGND VGND VPWR VPWR U$$1038/A sky130_fd_sc_hd__a22o_1
XU$$1048 U$$1048/A U$$1094/B VGND VGND VPWR VPWR U$$1048/X sky130_fd_sc_hd__xor2_1
XU$$1059 U$$98/B1 U$$1075/A2 U$$924/A1 U$$1075/B2 VGND VGND VPWR VPWR U$$1060/A sky130_fd_sc_hd__a22o_1
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1160 U$$3056/A1 VGND VGND VPWR VPWR U$$999/B1 sky130_fd_sc_hd__buf_4
Xfanout1171 U$$4424/A1 VGND VGND VPWR VPWR U$$4287/A1 sky130_fd_sc_hd__buf_6
XFILLER_78_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1182 U$$4011/A1 VGND VGND VPWR VPWR U$$38/A1 sky130_fd_sc_hd__buf_4
Xfanout1193 U$$1062/B VGND VGND VPWR VPWR U$$998/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_41_2 U$$2350/X U$$2483/X U$$2616/X VGND VGND VPWR VPWR dadda_fa_3_42_1/A
+ dadda_fa_3_41_3/A sky130_fd_sc_hd__fa_1
XFILLER_54_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_34_1 U$$740/X U$$873/X U$$1006/X VGND VGND VPWR VPWR dadda_fa_3_35_0/CIN
+ dadda_fa_3_34_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2250 U$$878/B1 U$$2252/A2 U$$745/A1 U$$2252/B2 VGND VGND VPWR VPWR U$$2251/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_11_0 U$$694/X input151/X dadda_fa_5_11_0/CIN VGND VGND VPWR VPWR dadda_fa_6_12_0/A
+ dadda_fa_6_11_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_27_0 U$$61/X U$$194/X U$$327/X VGND VGND VPWR VPWR dadda_fa_3_28_2/A dadda_fa_3_27_3/B
+ sky130_fd_sc_hd__fa_1
XU$$2261 U$$2261/A U$$2269/B VGND VGND VPWR VPWR U$$2261/X sky130_fd_sc_hd__xor2_1
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2272 U$$902/A1 U$$2272/A2 U$$902/B1 U$$2272/B2 VGND VGND VPWR VPWR U$$2273/A sky130_fd_sc_hd__a22o_1
XFILLER_90_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2283 U$$2283/A U$$2283/B VGND VGND VPWR VPWR U$$2283/X sky130_fd_sc_hd__xor2_1
XU$$2294 U$$922/B1 U$$2320/A2 U$$2707/A1 U$$2320/B2 VGND VGND VPWR VPWR U$$2295/A
+ sky130_fd_sc_hd__a22o_1
XU$$1560 U$$1560/A U$$1564/B VGND VGND VPWR VPWR U$$1560/X sky130_fd_sc_hd__xor2_1
XFILLER_50_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1571 U$$747/B1 U$$1587/A2 U$$749/B1 U$$1587/B2 VGND VGND VPWR VPWR U$$1572/A sky130_fd_sc_hd__a22o_1
XU$$1582 U$$1582/A U$$1584/B VGND VGND VPWR VPWR U$$1582/X sky130_fd_sc_hd__xor2_1
XFILLER_148_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1593 U$$632/B1 U$$1593/A2 U$$499/A1 U$$1593/B2 VGND VGND VPWR VPWR U$$1594/A sky130_fd_sc_hd__a22o_1
XFILLER_147_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1006 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_86_4 U$$3105/X U$$3238/X U$$3371/X VGND VGND VPWR VPWR dadda_fa_2_87_4/A
+ dadda_fa_2_86_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_79_3 U$$2293/X U$$2426/X U$$2559/X VGND VGND VPWR VPWR dadda_fa_2_80_1/B
+ dadda_fa_2_79_4/B sky130_fd_sc_hd__fa_1
XFILLER_98_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_56_2 dadda_fa_4_56_2/A dadda_fa_4_56_2/B dadda_fa_4_56_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_57_0/CIN dadda_fa_5_56_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$201 final_adder.U$$200/B final_adder.U$$971/B1 final_adder.U$$201/B1
+ VGND VGND VPWR VPWR final_adder.U$$201/X sky130_fd_sc_hd__a21o_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$212 final_adder.U$$212/A final_adder.U$$212/B VGND VGND VPWR VPWR
+ final_adder.U$$340/B sky130_fd_sc_hd__and2_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$223 final_adder.U$$222/B final_adder.U$$993/B1 final_adder.U$$223/B1
+ VGND VGND VPWR VPWR final_adder.U$$223/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_4_49_1 dadda_fa_4_49_1/A dadda_fa_4_49_1/B dadda_fa_4_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_50_0/B dadda_fa_5_49_1/B sky130_fd_sc_hd__fa_1
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$234 final_adder.U$$234/A final_adder.U$$234/B VGND VGND VPWR VPWR
+ final_adder.U$$362/B sky130_fd_sc_hd__and2_1
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$245 final_adder.U$$244/B final_adder.U$$245/A2 final_adder.U$$245/B1
+ VGND VGND VPWR VPWR final_adder.U$$245/X sky130_fd_sc_hd__a21o_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_26_0 dadda_fa_7_26_0/A dadda_fa_7_26_0/B dadda_fa_7_26_0/CIN VGND VGND
+ VPWR VPWR _323_/D _194_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$267 final_adder.U$$266/B final_adder.U$$141/X final_adder.U$$139/X
+ VGND VGND VPWR VPWR final_adder.U$$267/X sky130_fd_sc_hd__a21o_1
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$106 U$$654/A1 U$$120/A2 U$$654/B1 U$$120/B2 VGND VGND VPWR VPWR U$$107/A sky130_fd_sc_hd__a22o_1
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$278 final_adder.U$$280/B final_adder.U$$278/B VGND VGND VPWR VPWR
+ final_adder.U$$404/B sky130_fd_sc_hd__and2_1
XFILLER_85_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$117 U$$117/A U$$121/B VGND VGND VPWR VPWR U$$117/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$289 final_adder.U$$288/B final_adder.U$$163/X final_adder.U$$161/X
+ VGND VGND VPWR VPWR final_adder.U$$289/X sky130_fd_sc_hd__a21o_1
XU$$128 U$$539/A1 U$$98/A2 U$$539/B1 U$$98/B2 VGND VGND VPWR VPWR U$$129/A sky130_fd_sc_hd__a22o_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$139 U$$274/A VGND VGND VPWR VPWR U$$139/Y sky130_fd_sc_hd__inv_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_390_ _408_/CLK _390_/D VGND VGND VPWR VPWR _390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1024 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput230 c[76] VGND VGND VPWR VPWR input230/X sky130_fd_sc_hd__buf_2
Xdadda_fa_3_51_1 dadda_fa_3_51_1/A dadda_fa_3_51_1/B dadda_fa_3_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_0/CIN dadda_fa_4_51_2/A sky130_fd_sc_hd__fa_1
Xinput241 c[86] VGND VGND VPWR VPWR input241/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput252 c[96] VGND VGND VPWR VPWR input252/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_0_67_1 U$$540/X U$$673/X U$$806/X VGND VGND VPWR VPWR dadda_fa_1_68_5/CIN
+ dadda_fa_1_67_7/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_44_0 dadda_fa_3_44_0/A dadda_fa_3_44_0/B dadda_fa_3_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_0/B dadda_fa_4_44_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_36_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$790 final_adder.U$$790/A final_adder.U$$790/B VGND VGND VPWR VPWR
+ final_adder.U$$790/X sky130_fd_sc_hd__and2_1
XU$$640 U$$640/A1 U$$682/A2 U$$916/A1 U$$682/B2 VGND VGND VPWR VPWR U$$641/A sky130_fd_sc_hd__a22o_1
XFILLER_1_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$651 U$$651/A U$$651/B VGND VGND VPWR VPWR U$$651/X sky130_fd_sc_hd__xor2_1
XFILLER_16_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$662 U$$936/A1 U$$674/A2 U$$936/B1 U$$674/B2 VGND VGND VPWR VPWR U$$663/A sky130_fd_sc_hd__a22o_1
XU$$673 U$$673/A U$$685/A VGND VGND VPWR VPWR U$$673/X sky130_fd_sc_hd__xor2_1
XFILLER_72_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$684 U$$684/A VGND VGND VPWR VPWR U$$684/Y sky130_fd_sc_hd__inv_1
XU$$695 U$$8/B1 U$$743/A2 U$$697/A1 U$$743/B2 VGND VGND VPWR VPWR U$$696/A sky130_fd_sc_hd__a22o_1
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_101_0 dadda_fa_7_101_0/A dadda_fa_7_101_0/B dadda_fa_7_101_0/CIN VGND
+ VGND VPWR VPWR _398_/D _269_/D sky130_fd_sc_hd__fa_1
XFILLER_172_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_96_3 U$$3657/X U$$3790/X U$$3923/X VGND VGND VPWR VPWR dadda_fa_3_97_1/B
+ dadda_fa_3_96_3/B sky130_fd_sc_hd__fa_1
XFILLER_160_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_89_2 U$$4175/X U$$4308/X U$$4441/X VGND VGND VPWR VPWR dadda_fa_3_90_1/A
+ dadda_fa_3_89_3/A sky130_fd_sc_hd__fa_1
XU$$3285_1817 VGND VGND VPWR VPWR U$$3285_1817/HI U$$3285/B1 sky130_fd_sc_hd__conb_1
XFILLER_153_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_66_1 dadda_fa_5_66_1/A dadda_fa_5_66_1/B dadda_fa_5_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_67_0/B dadda_fa_7_66_0/A sky130_fd_sc_hd__fa_1
Xfanout408 U$$676/A2 VGND VGND VPWR VPWR U$$630/A2 sky130_fd_sc_hd__buf_4
Xfanout419 U$$4369/A2 VGND VGND VPWR VPWR U$$4373/A2 sky130_fd_sc_hd__buf_4
XFILLER_113_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_59_0 dadda_fa_5_59_0/A dadda_fa_5_59_0/B dadda_fa_5_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_60_0/A dadda_fa_6_59_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_58_8 dadda_fa_1_58_8/A dadda_fa_1_58_8/B dadda_fa_1_58_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_59_3/A dadda_fa_3_58_0/A sky130_fd_sc_hd__fa_2
XFILLER_67_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_105_0 U$$2876/Y U$$3010/X U$$3143/X VGND VGND VPWR VPWR dadda_fa_3_106_3/A
+ dadda_fa_3_105_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2080 U$$2080/A U$$2106/B VGND VGND VPWR VPWR U$$2080/X sky130_fd_sc_hd__xor2_1
XU$$2091 U$$995/A1 U$$2097/A2 U$$997/A1 U$$2097/B2 VGND VGND VPWR VPWR U$$2092/A sky130_fd_sc_hd__a22o_1
XFILLER_50_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1390 U$$2758/B1 U$$1426/A2 U$$2625/A1 U$$1426/B2 VGND VGND VPWR VPWR U$$1391/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_91_2 U$$2716/X U$$2849/X U$$2982/X VGND VGND VPWR VPWR dadda_fa_2_92_5/A
+ dadda_fa_3_91_0/A sky130_fd_sc_hd__fa_1
XFILLER_117_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_84_1 U$$1771/X U$$1904/X U$$2037/X VGND VGND VPWR VPWR dadda_fa_2_85_2/B
+ dadda_fa_2_84_4/B sky130_fd_sc_hd__fa_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_61_0 dadda_fa_4_61_0/A dadda_fa_4_61_0/B dadda_fa_4_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_62_0/A dadda_fa_5_61_1/A sky130_fd_sc_hd__fa_1
Xfanout920 U$$5/X VGND VGND VPWR VPWR U$$102/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout931 fanout938/X VGND VGND VPWR VPWR U$$3239/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_77_0 U$$1358/X U$$1491/X U$$1624/X VGND VGND VPWR VPWR dadda_fa_2_78_0/B
+ dadda_fa_2_77_3/B sky130_fd_sc_hd__fa_1
XFILLER_104_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout942 U$$4398/A1 VGND VGND VPWR VPWR U$$4259/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout953 U$$908/A1 VGND VGND VPWR VPWR U$$906/B1 sky130_fd_sc_hd__buf_6
Xfanout964 U$$4468/A1 VGND VGND VPWR VPWR U$$4331/A1 sky130_fd_sc_hd__buf_4
Xdadda_ha_2_104_2 U$$3540/X U$$3673/X VGND VGND VPWR VPWR dadda_fa_3_105_3/B dadda_fa_4_104_0/A
+ sky130_fd_sc_hd__ha_1
Xfanout975 input95/X VGND VGND VPWR VPWR fanout975/X sky130_fd_sc_hd__buf_6
Xfanout986 fanout993/X VGND VGND VPWR VPWR U$$487/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout997 fanout999/A VGND VGND VPWR VPWR U$$3775/A1 sky130_fd_sc_hd__buf_4
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3709 U$$3846/A1 U$$3791/A2 U$$3846/B1 U$$3791/B2 VGND VGND VPWR VPWR U$$3710/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_373_ _375_/CLK _373_/D VGND VGND VPWR VPWR _373_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_99_1 dadda_fa_3_99_1/A dadda_fa_3_99_1/B dadda_fa_3_99_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_100_0/CIN dadda_fa_4_99_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_76_0 dadda_fa_6_76_0/A dadda_fa_6_76_0/B dadda_fa_6_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_77_0/B dadda_fa_7_76_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$470 U$$470/A U$$504/B VGND VGND VPWR VPWR U$$470/X sky130_fd_sc_hd__xor2_1
XU$$481 U$$481/A1 U$$505/A2 U$$72/A1 U$$505/B2 VGND VGND VPWR VPWR U$$482/A sky130_fd_sc_hd__a22o_1
XU$$492 U$$492/A U$$498/B VGND VGND VPWR VPWR U$$492/X sky130_fd_sc_hd__xor2_1
XFILLER_149_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_94_0 U$$2722/X U$$2855/X U$$2988/X VGND VGND VPWR VPWR dadda_fa_3_95_0/B
+ dadda_fa_3_94_2/B sky130_fd_sc_hd__fa_1
XU$$4419_1857 VGND VGND VPWR VPWR U$$4419_1857/HI U$$4419/B sky130_fd_sc_hd__conb_1
Xdadda_fa_1_70_7 dadda_fa_1_70_7/A dadda_fa_1_70_7/B dadda_fa_1_70_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_71_2/CIN dadda_fa_2_70_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_63_6 dadda_fa_1_63_6/A dadda_fa_1_63_6/B dadda_fa_1_63_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_64_2/B dadda_fa_2_63_5/B sky130_fd_sc_hd__fa_1
XFILLER_86_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_56_5 U$$3178/X U$$3311/X U$$3444/X VGND VGND VPWR VPWR dadda_fa_2_57_2/A
+ dadda_fa_2_56_5/A sky130_fd_sc_hd__fa_1
XFILLER_83_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_49_4 U$$1701/X U$$1834/X U$$1967/X VGND VGND VPWR VPWR dadda_fa_2_50_2/A
+ dadda_fa_2_49_5/A sky130_fd_sc_hd__fa_1
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_19_2 dadda_fa_4_19_2/A dadda_fa_4_19_2/B dadda_ha_3_19_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_20_0/CIN dadda_fa_5_19_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_50_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_93_0 dadda_fa_7_93_0/A dadda_fa_7_93_0/B dadda_fa_7_93_0/CIN VGND VGND
+ VPWR VPWR _390_/D _261_/D sky130_fd_sc_hd__fa_2
XFILLER_137_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1704 fanout1708/X VGND VGND VPWR VPWR U$$517/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1715 fanout1718/X VGND VGND VPWR VPWR U$$4349/B1 sky130_fd_sc_hd__buf_4
XFILLER_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1726 input106/X VGND VGND VPWR VPWR U$$4486/A1 sky130_fd_sc_hd__buf_6
Xfanout1737 U$$370/B1 VGND VGND VPWR VPWR U$$3112/A1 sky130_fd_sc_hd__buf_2
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout750 U$$3439/B2 VGND VGND VPWR VPWR U$$3557/B2 sky130_fd_sc_hd__buf_4
Xfanout1748 U$$781/A1 VGND VGND VPWR VPWR U$$918/A1 sky130_fd_sc_hd__buf_6
Xfanout761 U$$3207/B2 VGND VGND VPWR VPWR U$$3199/B2 sky130_fd_sc_hd__buf_6
XU$$4207 U$$4207/A U$$4227/B VGND VGND VPWR VPWR U$$4207/X sky130_fd_sc_hd__xor2_1
Xfanout1759 U$$3382/A1 VGND VGND VPWR VPWR U$$4341/A1 sky130_fd_sc_hd__buf_2
Xfanout772 U$$3112/B2 VGND VGND VPWR VPWR U$$3108/B2 sky130_fd_sc_hd__buf_4
XU$$4218 U$$4353/B1 U$$4240/A2 U$$4220/A1 U$$4240/B2 VGND VGND VPWR VPWR U$$4219/A
+ sky130_fd_sc_hd__a22o_1
Xfanout783 U$$2882/X VGND VGND VPWR VPWR U$$2991/B2 sky130_fd_sc_hd__buf_6
XU$$4229 U$$4229/A U$$4231/B VGND VGND VPWR VPWR U$$4229/X sky130_fd_sc_hd__xor2_1
XFILLER_58_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout794 U$$386/B2 VGND VGND VPWR VPWR U$$338/B2 sky130_fd_sc_hd__buf_2
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3506 U$$3506/A U$$3506/B VGND VGND VPWR VPWR U$$3506/X sky130_fd_sc_hd__xor2_1
XFILLER_19_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3517 U$$4476/A1 U$$3557/A2 U$$4478/A1 U$$3557/B2 VGND VGND VPWR VPWR U$$3518/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3528 U$$3528/A U$$3548/B VGND VGND VPWR VPWR U$$3528/X sky130_fd_sc_hd__xor2_1
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3539 U$$4359/B1 U$$3549/A2 U$$4226/A1 U$$3549/B2 VGND VGND VPWR VPWR U$$3540/A
+ sky130_fd_sc_hd__a22o_1
XU$$2805 U$$2805/A U$$2805/B VGND VGND VPWR VPWR U$$2805/X sky130_fd_sc_hd__xor2_1
XFILLER_74_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2816 U$$4049/A1 U$$2872/A2 U$$4460/B1 U$$2872/B2 VGND VGND VPWR VPWR U$$2817/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2827 U$$2827/A U$$2841/B VGND VGND VPWR VPWR U$$2827/X sky130_fd_sc_hd__xor2_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2838 U$$2973/B1 U$$2840/A2 U$$2840/A1 U$$2840/B2 VGND VGND VPWR VPWR U$$2839/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2849 U$$2849/A U$$2876/A VGND VGND VPWR VPWR U$$2849/X sky130_fd_sc_hd__xor2_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_21_2 U$$847/X U$$980/X U$$1113/X VGND VGND VPWR VPWR dadda_fa_4_22_1/A
+ dadda_fa_4_21_2/B sky130_fd_sc_hd__fa_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_356_ _356_/CLK _356_/D VGND VGND VPWR VPWR _356_/Q sky130_fd_sc_hd__dfxtp_1
X_287_ _415_/CLK _287_/D VGND VGND VPWR VPWR _287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_73_5 dadda_fa_2_73_5/A dadda_fa_2_73_5/B dadda_fa_2_73_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_2/A dadda_fa_4_73_0/A sky130_fd_sc_hd__fa_1
XFILLER_111_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_66_4 dadda_fa_2_66_4/A dadda_fa_2_66_4/B dadda_fa_2_66_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_1/CIN dadda_fa_3_66_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_59_3 dadda_fa_2_59_3/A dadda_fa_2_59_3/B dadda_fa_2_59_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_1/B dadda_fa_3_59_3/B sky130_fd_sc_hd__fa_1
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 a[13] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_29_1 dadda_fa_5_29_1/A dadda_fa_5_29_1/B dadda_fa_5_29_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_30_0/B dadda_fa_7_29_0/A sky130_fd_sc_hd__fa_1
XFILLER_51_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$3 _299_/Q _171_/Q VGND VGND VPWR VPWR final_adder.U$$3/COUT final_adder.U$$3/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_173_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_103_1 dadda_fa_5_103_1/A dadda_fa_5_103_1/B dadda_fa_5_103_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_104_0/B dadda_fa_7_103_0/A sky130_fd_sc_hd__fa_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput320 output320/A VGND VGND VPWR VPWR o[41] sky130_fd_sc_hd__buf_2
Xoutput331 output331/A VGND VGND VPWR VPWR o[51] sky130_fd_sc_hd__buf_2
XFILLER_126_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput342 output342/A VGND VGND VPWR VPWR o[61] sky130_fd_sc_hd__buf_2
XFILLER_161_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput353 output353/A VGND VGND VPWR VPWR o[71] sky130_fd_sc_hd__buf_2
Xoutput364 output364/A VGND VGND VPWR VPWR o[81] sky130_fd_sc_hd__buf_2
Xoutput375 output375/A VGND VGND VPWR VPWR o[91] sky130_fd_sc_hd__buf_2
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_3 U$$3188/X U$$3321/X U$$3454/X VGND VGND VPWR VPWR dadda_fa_2_62_1/B
+ dadda_fa_2_61_4/B sky130_fd_sc_hd__fa_1
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_54_2 U$$1578/X U$$1711/X U$$1844/X VGND VGND VPWR VPWR dadda_fa_2_55_1/A
+ dadda_fa_2_54_4/A sky130_fd_sc_hd__fa_1
XFILLER_56_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_31_1 dadda_fa_4_31_1/A dadda_fa_4_31_1/B dadda_fa_4_31_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_32_0/B dadda_fa_5_31_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_47_1 U$$500/X U$$633/X U$$766/X VGND VGND VPWR VPWR dadda_fa_2_48_1/CIN
+ dadda_fa_2_47_4/B sky130_fd_sc_hd__fa_1
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_24_0 dadda_fa_4_24_0/A dadda_fa_4_24_0/B dadda_fa_4_24_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_25_0/A dadda_fa_5_24_1/A sky130_fd_sc_hd__fa_1
XFILLER_70_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_210_ _344_/CLK _210_/D VGND VGND VPWR VPWR _210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$280_1810 VGND VGND VPWR VPWR U$$280_1810/HI U$$280/A1 sky130_fd_sc_hd__conb_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4107_1831 VGND VGND VPWR VPWR U$$4107_1831/HI U$$4107/B1 sky130_fd_sc_hd__conb_1
XFILLER_168_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_76_3 dadda_fa_3_76_3/A dadda_fa_3_76_3/B dadda_fa_3_76_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_1/B dadda_fa_4_76_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1501 input14/X VGND VGND VPWR VPWR U$$1455/B sky130_fd_sc_hd__buf_4
Xdadda_fa_3_69_2 dadda_fa_3_69_2/A dadda_fa_3_69_2/B dadda_fa_3_69_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_1/A dadda_fa_4_69_2/B sky130_fd_sc_hd__fa_1
Xfanout1512 U$$4410/A1 VGND VGND VPWR VPWR U$$3314/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1523 U$$2897/B1 VGND VGND VPWR VPWR U$$2625/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1534 input125/X VGND VGND VPWR VPWR U$$4404/A1 sky130_fd_sc_hd__buf_6
XFILLER_120_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1545 U$$3559/A1 VGND VGND VPWR VPWR U$$3285/A1 sky130_fd_sc_hd__buf_4
Xfanout1556 U$$4514/A1 VGND VGND VPWR VPWR U$$539/B1 sky130_fd_sc_hd__buf_4
XU$$4004 U$$4004/A U$$4006/B VGND VGND VPWR VPWR U$$4004/X sky130_fd_sc_hd__xor2_1
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1567 U$$4512/A1 VGND VGND VPWR VPWR U$$2183/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4015 U$$4152/A1 U$$4105/A2 U$$4152/B1 U$$4105/B2 VGND VGND VPWR VPWR U$$4016/A
+ sky130_fd_sc_hd__a22o_1
XU$$4026 U$$4026/A U$$4026/B VGND VGND VPWR VPWR U$$4026/X sky130_fd_sc_hd__xor2_1
Xfanout580 U$$2147/A2 VGND VGND VPWR VPWR U$$2107/A2 sky130_fd_sc_hd__buf_6
Xfanout1578 U$$566/A1 VGND VGND VPWR VPWR U$$18/A1 sky130_fd_sc_hd__clkbuf_4
XU$$4037 U$$4174/A1 U$$4045/A2 U$$4176/A1 U$$4045/B2 VGND VGND VPWR VPWR U$$4038/A
+ sky130_fd_sc_hd__a22o_1
Xfanout591 U$$2052/A2 VGND VGND VPWR VPWR U$$2044/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout1589 U$$77/B VGND VGND VPWR VPWR U$$81/B sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_6_39_0 dadda_fa_6_39_0/A dadda_fa_6_39_0/B dadda_fa_6_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_40_0/B dadda_fa_7_39_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4048 U$$4048/A U$$4098/B VGND VGND VPWR VPWR U$$4048/X sky130_fd_sc_hd__xor2_1
XU$$3303 U$$3303/A U$$3349/B VGND VGND VPWR VPWR U$$3303/X sky130_fd_sc_hd__xor2_1
XU$$3314 U$$3314/A1 U$$3390/A2 U$$3314/B1 U$$3390/B2 VGND VGND VPWR VPWR U$$3315/A
+ sky130_fd_sc_hd__a22o_1
XU$$4059 U$$4196/A1 U$$4081/A2 U$$4196/B1 U$$4081/B2 VGND VGND VPWR VPWR U$$4060/A
+ sky130_fd_sc_hd__a22o_1
XU$$3325 U$$3325/A U$$3335/B VGND VGND VPWR VPWR U$$3325/X sky130_fd_sc_hd__xor2_1
XFILLER_47_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3336 U$$4158/A1 U$$3340/A2 U$$4295/B1 U$$3340/B2 VGND VGND VPWR VPWR U$$3337/A
+ sky130_fd_sc_hd__a22o_1
XU$$2602 U$$2602/A VGND VGND VPWR VPWR U$$2602/Y sky130_fd_sc_hd__inv_1
XU$$3347 U$$3347/A U$$3391/B VGND VGND VPWR VPWR U$$3347/X sky130_fd_sc_hd__xor2_1
XU$$3358 U$$3630/B1 U$$3372/A2 U$$3495/B1 U$$3372/B2 VGND VGND VPWR VPWR U$$3359/A
+ sky130_fd_sc_hd__a22o_1
XU$$2613 U$$4257/A1 U$$2667/A2 U$$3298/B1 U$$2667/B2 VGND VGND VPWR VPWR U$$2614/A
+ sky130_fd_sc_hd__a22o_1
XU$$3369 U$$3369/A U$$3373/B VGND VGND VPWR VPWR U$$3369/X sky130_fd_sc_hd__xor2_1
XU$$2624 U$$2624/A U$$2662/B VGND VGND VPWR VPWR U$$2624/X sky130_fd_sc_hd__xor2_1
XFILLER_61_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2635 U$$3181/B1 U$$2681/A2 U$$32/B1 U$$2681/B2 VGND VGND VPWR VPWR U$$2636/A sky130_fd_sc_hd__a22o_1
XU$$1901 U$$942/A1 U$$1911/A2 U$$2175/B1 U$$1911/B2 VGND VGND VPWR VPWR U$$1902/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2646 U$$2646/A U$$2724/B VGND VGND VPWR VPWR U$$2646/X sky130_fd_sc_hd__xor2_1
XU$$1912 U$$1912/A U$$1918/A VGND VGND VPWR VPWR U$$1912/X sky130_fd_sc_hd__xor2_1
XU$$2657 U$$602/A1 U$$2665/A2 U$$3205/B1 U$$2665/B2 VGND VGND VPWR VPWR U$$2658/A
+ sky130_fd_sc_hd__a22o_1
XU$$1923 U$$1921/B U$$1918/A input21/X U$$1918/Y VGND VGND VPWR VPWR U$$1923/X sky130_fd_sc_hd__a22o_1
XU$$2668 U$$2668/A U$$2668/B VGND VGND VPWR VPWR U$$2668/X sky130_fd_sc_hd__xor2_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1934 U$$973/B1 U$$1980/A2 U$$840/A1 U$$1980/B2 VGND VGND VPWR VPWR U$$1935/A sky130_fd_sc_hd__a22o_1
XU$$2679 U$$76/A1 U$$2679/A2 U$$78/A1 U$$2679/B2 VGND VGND VPWR VPWR U$$2680/A sky130_fd_sc_hd__a22o_1
XU$$1945 U$$1945/A U$$1971/B VGND VGND VPWR VPWR U$$1945/X sky130_fd_sc_hd__xor2_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1956 U$$997/A1 U$$1964/A2 U$$997/B1 U$$1964/B2 VGND VGND VPWR VPWR U$$1957/A sky130_fd_sc_hd__a22o_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1967 U$$1967/A U$$1971/B VGND VGND VPWR VPWR U$$1967/X sky130_fd_sc_hd__xor2_1
XU$$1978 U$$745/A1 U$$2014/A2 U$$745/B1 U$$2014/B2 VGND VGND VPWR VPWR U$$1979/A sky130_fd_sc_hd__a22o_1
X_408_ _408_/CLK _408_/D VGND VGND VPWR VPWR _408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1989 U$$1989/A U$$2007/B VGND VGND VPWR VPWR U$$1989/X sky130_fd_sc_hd__xor2_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_339_ _353_/CLK _339_/D VGND VGND VPWR VPWR _339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_948 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_71_2 dadda_fa_2_71_2/A dadda_fa_2_71_2/B dadda_fa_2_71_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_1/A dadda_fa_3_71_3/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_64_1 dadda_fa_2_64_1/A dadda_fa_2_64_1/B dadda_fa_2_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_0/CIN dadda_fa_3_64_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$608 final_adder.U$$616/B final_adder.U$$608/B VGND VGND VPWR VPWR
+ final_adder.U$$712/A sky130_fd_sc_hd__and2_1
XFILLER_110_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$619 final_adder.U$$610/A final_adder.U$$503/X final_adder.U$$495/X
+ VGND VGND VPWR VPWR final_adder.U$$619/X sky130_fd_sc_hd__a21o_2
XFILLER_57_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_41_0 dadda_fa_5_41_0/A dadda_fa_5_41_0/B dadda_fa_5_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_42_0/A dadda_fa_6_41_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_57_0 dadda_fa_2_57_0/A dadda_fa_2_57_0/B dadda_fa_2_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_0/B dadda_fa_3_57_2/B sky130_fd_sc_hd__fa_1
XU$$30 U$$30/A1 U$$80/A2 U$$32/A1 U$$80/B2 VGND VGND VPWR VPWR U$$31/A sky130_fd_sc_hd__a22o_1
XU$$41 U$$41/A U$$77/B VGND VGND VPWR VPWR U$$41/X sky130_fd_sc_hd__xor2_1
XU$$52 U$$52/A1 U$$86/A2 U$$54/A1 U$$86/B2 VGND VGND VPWR VPWR U$$53/A sky130_fd_sc_hd__a22o_1
XU$$63 U$$63/A U$$97/B VGND VGND VPWR VPWR U$$63/X sky130_fd_sc_hd__xor2_1
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$74 U$$74/A1 U$$74/A2 U$$74/B1 U$$74/B2 VGND VGND VPWR VPWR U$$75/A sky130_fd_sc_hd__a22o_1
XU$$3870 U$$3870/A1 U$$3872/A2 U$$3870/B1 U$$3872/B2 VGND VGND VPWR VPWR U$$3871/A
+ sky130_fd_sc_hd__a22o_1
XU$$85 U$$85/A U$$87/B VGND VGND VPWR VPWR U$$85/X sky130_fd_sc_hd__xor2_1
XU$$96 U$$96/A1 U$$96/A2 U$$98/A1 U$$96/B2 VGND VGND VPWR VPWR U$$97/A sky130_fd_sc_hd__a22o_1
XU$$3881 U$$3881/A U$$3925/B VGND VGND VPWR VPWR U$$3881/X sky130_fd_sc_hd__xor2_1
XU$$3892 U$$4027/B1 U$$3892/A2 U$$4442/A1 U$$3892/B2 VGND VGND VPWR VPWR U$$3893/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4503_1899 VGND VGND VPWR VPWR U$$4503_1899/HI U$$4503/B sky130_fd_sc_hd__conb_1
XFILLER_122_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_86_2 dadda_fa_4_86_2/A dadda_fa_4_86_2/B dadda_fa_4_86_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_87_0/CIN dadda_fa_5_86_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_79_1 dadda_fa_4_79_1/A dadda_fa_4_79_1/B dadda_fa_4_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_80_0/B dadda_fa_5_79_1/B sky130_fd_sc_hd__fa_1
XFILLER_133_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3011_1813 VGND VGND VPWR VPWR U$$3011_1813/HI U$$3011/B1 sky130_fd_sc_hd__conb_1
Xdadda_fa_7_56_0 dadda_fa_7_56_0/A dadda_fa_7_56_0/B dadda_fa_7_56_0/CIN VGND VGND
+ VPWR VPWR _353_/D _224_/D sky130_fd_sc_hd__fa_1
XFILLER_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1208 U$$2578/A1 U$$1230/A2 U$$388/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1209/A
+ sky130_fd_sc_hd__a22o_1
XU$$1219 U$$1219/A U$$1221/B VGND VGND VPWR VPWR U$$1219/X sky130_fd_sc_hd__xor2_1
XFILLER_44_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_815 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1013 final_adder.U$$242/A final_adder.U$$623/X final_adder.U$$243/A2
+ VGND VGND VPWR VPWR final_adder.U$$1037/B sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$1024 final_adder.U$$0/SUM final_adder.U$$1024/B VGND VGND VPWR VPWR
+ output257/A sky130_fd_sc_hd__xor2_1
XFILLER_8_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1035 final_adder.U$$244/B final_adder.U$$1035/B VGND VGND VPWR VPWR
+ output279/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1046 final_adder.U$$232/A final_adder.U$$733/X VGND VGND VPWR VPWR
+ output299/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1057 final_adder.U$$222/B final_adder.U$$993/X VGND VGND VPWR VPWR
+ output311/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1068 final_adder.U$$210/A final_adder.U$$823/X VGND VGND VPWR VPWR
+ output323/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1079 final_adder.U$$200/B final_adder.U$$971/X VGND VGND VPWR VPWR
+ output335/A sky130_fd_sc_hd__xor2_1
XFILLER_124_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_81_1 dadda_fa_3_81_1/A dadda_fa_3_81_1/B dadda_fa_3_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_0/CIN dadda_fa_4_81_2/A sky130_fd_sc_hd__fa_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_74_0 dadda_fa_3_74_0/A dadda_fa_3_74_0/B dadda_fa_3_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_0/B dadda_fa_4_74_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1320 U$$955/B VGND VGND VPWR VPWR U$$925/B sky130_fd_sc_hd__buf_8
XFILLER_87_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1331 input49/X VGND VGND VPWR VPWR U$$3607/B sky130_fd_sc_hd__buf_6
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1342 U$$3561/A VGND VGND VPWR VPWR U$$3558/B sky130_fd_sc_hd__buf_6
XFILLER_93_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1353 U$$3391/B VGND VGND VPWR VPWR U$$3424/A sky130_fd_sc_hd__buf_6
Xfanout1364 input42/X VGND VGND VPWR VPWR fanout1364/X sky130_fd_sc_hd__buf_6
XFILLER_78_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1010 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1375 input38/X VGND VGND VPWR VPWR U$$2938/B sky130_fd_sc_hd__buf_6
XFILLER_94_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1386 fanout1391/X VGND VGND VPWR VPWR U$$2877/A sky130_fd_sc_hd__buf_6
XU$$3100 U$$3372/B1 U$$3108/A2 U$$3239/A1 U$$3108/B2 VGND VGND VPWR VPWR U$$3101/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1397 U$$182/B VGND VGND VPWR VPWR U$$180/B sky130_fd_sc_hd__buf_4
XU$$3111 U$$3111/A U$$3151/A VGND VGND VPWR VPWR U$$3111/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_110_1 dadda_fa_4_110_1/A dadda_fa_4_110_1/B dadda_fa_4_110_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_111_0/B dadda_fa_5_110_1/B sky130_fd_sc_hd__fa_1
XU$$3122 U$$517/B1 U$$3122/A2 U$$384/A1 U$$3122/B2 VGND VGND VPWR VPWR U$$3123/A sky130_fd_sc_hd__a22o_1
XU$$3133 U$$3133/A U$$3150/A VGND VGND VPWR VPWR U$$3133/X sky130_fd_sc_hd__xor2_1
XU$$3144 U$$3418/A1 U$$3144/A2 U$$3418/B1 U$$3144/B2 VGND VGND VPWR VPWR U$$3145/A
+ sky130_fd_sc_hd__a22o_1
XU$$3155 U$$3153/Y input41/X U$$3151/A U$$3154/X U$$3151/Y VGND VGND VPWR VPWR U$$3155/X
+ sky130_fd_sc_hd__a32o_2
XU$$2410 U$$2410/A U$$2456/B VGND VGND VPWR VPWR U$$2410/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_36_5 input186/X dadda_fa_2_36_5/B dadda_fa_2_36_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_37_2/A dadda_fa_4_36_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_103_0 dadda_fa_4_103_0/A dadda_fa_4_103_0/B dadda_fa_4_103_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_104_0/A dadda_fa_5_103_1/A sky130_fd_sc_hd__fa_1
XU$$3166 U$$3166/A U$$3210/B VGND VGND VPWR VPWR U$$3166/X sky130_fd_sc_hd__xor2_1
XU$$2421 U$$4476/A1 U$$2463/A2 U$$4478/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2422/A
+ sky130_fd_sc_hd__a22o_1
XU$$2432 U$$2432/A U$$2466/A VGND VGND VPWR VPWR U$$2432/X sky130_fd_sc_hd__xor2_1
XFILLER_62_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3177 U$$4410/A1 U$$3255/A2 U$$4412/A1 U$$3255/B2 VGND VGND VPWR VPWR U$$3178/A
+ sky130_fd_sc_hd__a22o_1
XU$$3188 U$$3188/A U$$3196/B VGND VGND VPWR VPWR U$$3188/X sky130_fd_sc_hd__xor2_1
XU$$2443 U$$2578/B1 U$$2443/A2 U$$2443/B1 U$$2443/B2 VGND VGND VPWR VPWR U$$2444/A
+ sky130_fd_sc_hd__a22o_1
XU$$2454 U$$2454/A U$$2456/B VGND VGND VPWR VPWR U$$2454/X sky130_fd_sc_hd__xor2_1
XU$$3199 U$$4158/A1 U$$3199/A2 U$$4295/B1 U$$3199/B2 VGND VGND VPWR VPWR U$$3200/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1720 U$$74/B1 U$$1720/A2 U$$215/A1 U$$1720/B2 VGND VGND VPWR VPWR U$$1721/A sky130_fd_sc_hd__a22o_1
XU$$2465 U$$2465/A VGND VGND VPWR VPWR U$$2465/Y sky130_fd_sc_hd__inv_1
XU$$1731 U$$1731/A U$$1741/B VGND VGND VPWR VPWR U$$1731/X sky130_fd_sc_hd__xor2_1
XU$$2476 U$$3846/A1 U$$2546/A2 U$$971/A1 U$$2546/B2 VGND VGND VPWR VPWR U$$2477/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2487 U$$2487/A U$$2529/B VGND VGND VPWR VPWR U$$2487/X sky130_fd_sc_hd__xor2_1
XU$$1742 U$$3249/A1 U$$1758/A2 U$$920/B1 U$$1758/B2 VGND VGND VPWR VPWR U$$1743/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2498 U$$852/B1 U$$2540/A2 U$$854/B1 U$$2540/B2 VGND VGND VPWR VPWR U$$2499/A sky130_fd_sc_hd__a22o_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1753 U$$1753/A U$$1761/B VGND VGND VPWR VPWR U$$1753/X sky130_fd_sc_hd__xor2_1
XU$$1764 U$$805/A1 U$$1778/A2 U$$805/B1 U$$1778/B2 VGND VGND VPWR VPWR U$$1765/A sky130_fd_sc_hd__a22o_1
XU$$1775 U$$1775/A U$$1777/B VGND VGND VPWR VPWR U$$1775/X sky130_fd_sc_hd__xor2_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1786 U$$1784/B U$$1741/B input19/X U$$1781/Y VGND VGND VPWR VPWR U$$1786/X sky130_fd_sc_hd__a22o_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1797 U$$3030/A1 U$$1831/A2 U$$3030/B1 U$$1831/B2 VGND VGND VPWR VPWR U$$1798/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_96_1 dadda_fa_5_96_1/A dadda_fa_5_96_1/B dadda_fa_5_96_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_97_0/B dadda_fa_7_96_0/A sky130_fd_sc_hd__fa_1
Xinput30 a[36] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput41 a[46] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_1
Xinput52 a[56] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_1
Xinput63 a[8] VGND VGND VPWR VPWR U$$549/A sky130_fd_sc_hd__buf_2
XFILLER_128_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_89_0 dadda_fa_5_89_0/A dadda_fa_5_89_0/B dadda_fa_5_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_90_0/A dadda_fa_6_89_0/CIN sky130_fd_sc_hd__fa_1
Xinput74 b[18] VGND VGND VPWR VPWR input74/X sky130_fd_sc_hd__buf_2
Xinput85 b[28] VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__buf_6
Xinput96 b[38] VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$405 final_adder.U$$404/B final_adder.U$$283/X final_adder.U$$279/X
+ VGND VGND VPWR VPWR final_adder.U$$405/X sky130_fd_sc_hd__a21o_1
XFILLER_111_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$416 final_adder.U$$420/B final_adder.U$$416/B VGND VGND VPWR VPWR
+ final_adder.U$$540/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$427 final_adder.U$$426/B final_adder.U$$305/X final_adder.U$$301/X
+ VGND VGND VPWR VPWR final_adder.U$$427/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$438 final_adder.U$$442/B final_adder.U$$438/B VGND VGND VPWR VPWR
+ final_adder.U$$562/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$449 final_adder.U$$448/B final_adder.U$$327/X final_adder.U$$323/X
+ VGND VGND VPWR VPWR final_adder.U$$449/X sky130_fd_sc_hd__a21o_1
XFILLER_38_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4390 U$$4390/A1 U$$4388/X U$$4392/A1 U$$4428/B2 VGND VGND VPWR VPWR U$$4391/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2609_1806 VGND VGND VPWR VPWR U$$2609_1806/HI U$$2609/A1 sky130_fd_sc_hd__conb_1
XFILLER_25_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_91_0 dadda_fa_4_91_0/A dadda_fa_4_91_0/B dadda_fa_4_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_92_0/A dadda_fa_5_91_1/A sky130_fd_sc_hd__fa_1
XFILLER_148_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_105_2 U$$4473/X input135/X dadda_fa_3_105_2/CIN VGND VGND VPWR VPWR dadda_fa_4_106_1/A
+ dadda_fa_4_105_2/B sky130_fd_sc_hd__fa_1
XFILLER_164_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_119_0 dadda_fa_6_119_0/A dadda_fa_6_119_0/B dadda_fa_6_119_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_120_0/B dadda_fa_7_119_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_169_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$961 final_adder.U$$190/A final_adder.U$$803/X final_adder.U$$961/B1
+ VGND VGND VPWR VPWR final_adder.U$$961/X sky130_fd_sc_hd__a21o_1
XFILLER_17_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$800 U$$800/A U$$804/B VGND VGND VPWR VPWR U$$800/X sky130_fd_sc_hd__xor2_1
XFILLER_29_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$811 U$$811/A1 U$$817/A2 U$$811/B1 U$$817/B2 VGND VGND VPWR VPWR U$$812/A sky130_fd_sc_hd__a22o_1
XFILLER_91_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$983 final_adder.U$$212/A final_adder.U$$825/X final_adder.U$$983/B1
+ VGND VGND VPWR VPWR final_adder.U$$983/X sky130_fd_sc_hd__a21o_1
XFILLER_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$822 U$$822/A VGND VGND VPWR VPWR U$$822/Y sky130_fd_sc_hd__inv_1
XFILLER_16_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_39_3 dadda_fa_3_39_3/A dadda_fa_3_39_3/B dadda_fa_3_39_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_1/B dadda_fa_4_39_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$833 U$$833/A U$$875/B VGND VGND VPWR VPWR U$$833/X sky130_fd_sc_hd__xor2_1
XFILLER_17_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$844 U$$22/A1 U$$876/A2 U$$24/A1 U$$876/B2 VGND VGND VPWR VPWR U$$845/A sky130_fd_sc_hd__a22o_1
XU$$855 U$$855/A U$$925/B VGND VGND VPWR VPWR U$$855/X sky130_fd_sc_hd__xor2_1
XU$$866 U$$866/A1 U$$902/A2 U$$868/A1 U$$902/B2 VGND VGND VPWR VPWR U$$867/A sky130_fd_sc_hd__a22o_1
XFILLER_44_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1005 U$$46/A1 U$$979/A2 U$$48/A1 U$$979/B2 VGND VGND VPWR VPWR U$$1006/A sky130_fd_sc_hd__a22o_1
XFILLER_32_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1016 U$$1016/A U$$982/B VGND VGND VPWR VPWR U$$1016/X sky130_fd_sc_hd__xor2_1
XU$$877 U$$877/A U$$913/B VGND VGND VPWR VPWR U$$877/X sky130_fd_sc_hd__xor2_1
XU$$1027 U$$66/B1 U$$997/A2 U$$892/A1 U$$997/B2 VGND VGND VPWR VPWR U$$1028/A sky130_fd_sc_hd__a22o_1
XU$$888 U$$64/B1 U$$898/A2 U$$66/B1 U$$898/B2 VGND VGND VPWR VPWR U$$889/A sky130_fd_sc_hd__a22o_1
XU$$899 U$$899/A U$$925/B VGND VGND VPWR VPWR U$$899/X sky130_fd_sc_hd__xor2_1
XFILLER_73_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1038 U$$1038/A U$$982/B VGND VGND VPWR VPWR U$$1038/X sky130_fd_sc_hd__xor2_1
XU$$1049 U$$773/B1 U$$1087/A2 U$$640/A1 U$$1087/B2 VGND VGND VPWR VPWR U$$1050/A sky130_fd_sc_hd__a22o_1
XFILLER_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1150 U$$3056/B1 VGND VGND VPWR VPWR U$$864/B1 sky130_fd_sc_hd__clkbuf_4
Xdadda_ha_2_28_3 U$$1260/X U$$1393/X VGND VGND VPWR VPWR dadda_fa_3_29_2/CIN dadda_fa_4_28_0/A
+ sky130_fd_sc_hd__ha_1
Xfanout1161 U$$4424/B1 VGND VGND VPWR VPWR U$$3056/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1172 U$$40/A1 VGND VGND VPWR VPWR U$$314/A1 sky130_fd_sc_hd__buf_4
Xfanout1183 U$$4422/A1 VGND VGND VPWR VPWR U$$4011/A1 sky130_fd_sc_hd__buf_6
Xfanout1194 U$$990/B VGND VGND VPWR VPWR U$$1062/B sky130_fd_sc_hd__buf_6
XFILLER_82_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_41_3 U$$2749/X input192/X dadda_fa_2_41_3/CIN VGND VGND VPWR VPWR dadda_fa_3_42_1/B
+ dadda_fa_3_41_3/B sky130_fd_sc_hd__fa_1
XFILLER_82_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_34_2 U$$1139/X U$$1272/X U$$1405/X VGND VGND VPWR VPWR dadda_fa_3_35_1/A
+ dadda_fa_3_34_3/A sky130_fd_sc_hd__fa_1
XU$$2240 U$$870/A1 U$$2252/A2 U$$50/A1 U$$2252/B2 VGND VGND VPWR VPWR U$$2241/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_11_1 dadda_fa_5_11_1/A dadda_fa_5_11_1/B dadda_ha_4_11_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_12_0/B dadda_fa_7_11_0/A sky130_fd_sc_hd__fa_1
XU$$2251 U$$2251/A U$$2253/B VGND VGND VPWR VPWR U$$2251/X sky130_fd_sc_hd__xor2_1
XFILLER_35_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2262 U$$70/A1 U$$2272/A2 U$$70/B1 U$$2272/B2 VGND VGND VPWR VPWR U$$2263/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_27_1 U$$460/X U$$593/X U$$726/X VGND VGND VPWR VPWR dadda_fa_3_28_2/B
+ dadda_fa_3_27_3/CIN sky130_fd_sc_hd__fa_1
XU$$2273 U$$2273/A U$$2273/B VGND VGND VPWR VPWR U$$2273/X sky130_fd_sc_hd__xor2_1
XU$$2284 U$$3515/B1 U$$2326/A2 U$$3382/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2285/A
+ sky130_fd_sc_hd__a22o_1
XU$$2295 U$$2295/A U$$2301/B VGND VGND VPWR VPWR U$$2295/X sky130_fd_sc_hd__xor2_1
XU$$1550 U$$1550/A U$$1568/B VGND VGND VPWR VPWR U$$1550/X sky130_fd_sc_hd__xor2_1
XU$$1561 U$$465/A1 U$$1563/A2 U$$56/A1 U$$1563/B2 VGND VGND VPWR VPWR U$$1562/A sky130_fd_sc_hd__a22o_1
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1572 U$$1572/A U$$1584/B VGND VGND VPWR VPWR U$$1572/X sky130_fd_sc_hd__xor2_1
XFILLER_22_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1583 U$$76/A1 U$$1587/A2 U$$78/A1 U$$1587/B2 VGND VGND VPWR VPWR U$$1584/A sky130_fd_sc_hd__a22o_1
XU$$1594 U$$1594/A U$$1594/B VGND VGND VPWR VPWR U$$1594/X sky130_fd_sc_hd__xor2_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_79_4 U$$2692/X U$$2825/X U$$2958/X VGND VGND VPWR VPWR dadda_fa_2_80_1/CIN
+ dadda_fa_2_79_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$202 final_adder.U$$202/A final_adder.U$$202/B VGND VGND VPWR VPWR
+ final_adder.U$$330/B sky130_fd_sc_hd__and2_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$213 final_adder.U$$212/B final_adder.U$$983/B1 final_adder.U$$213/B1
+ VGND VGND VPWR VPWR final_adder.U$$213/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$224 final_adder.U$$224/A final_adder.U$$224/B VGND VGND VPWR VPWR
+ final_adder.U$$352/B sky130_fd_sc_hd__and2_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_49_2 dadda_fa_4_49_2/A dadda_fa_4_49_2/B dadda_fa_4_49_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_50_0/CIN dadda_fa_5_49_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$235 final_adder.U$$234/B final_adder.U$$235/A2 final_adder.U$$235/B1
+ VGND VGND VPWR VPWR final_adder.U$$235/X sky130_fd_sc_hd__a21o_1
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$246 final_adder.U$$8/SUM final_adder.U$$9/SUM VGND VGND VPWR VPWR
+ final_adder.U$$374/B sky130_fd_sc_hd__and2_1
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$268 final_adder.U$$270/B final_adder.U$$268/B VGND VGND VPWR VPWR
+ final_adder.U$$394/B sky130_fd_sc_hd__and2_1
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$107 U$$107/A U$$121/B VGND VGND VPWR VPWR U$$107/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$279 final_adder.U$$278/B final_adder.U$$153/X final_adder.U$$151/X
+ VGND VGND VPWR VPWR final_adder.U$$279/X sky130_fd_sc_hd__a21o_1
XFILLER_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$118 U$$253/B1 U$$120/A2 U$$120/A1 U$$120/B2 VGND VGND VPWR VPWR U$$119/A sky130_fd_sc_hd__a22o_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$129 U$$129/A U$$99/B VGND VGND VPWR VPWR U$$129/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_19_0 dadda_fa_7_19_0/A dadda_fa_7_19_0/B dadda_fa_7_19_0/CIN VGND VGND
+ VPWR VPWR _316_/D _187_/D sky130_fd_sc_hd__fa_2
XFILLER_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1032 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_110_0 dadda_fa_3_110_0/A U$$3286/X U$$3419/X VGND VGND VPWR VPWR dadda_fa_4_111_0/CIN
+ dadda_fa_4_110_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1787_1794 VGND VGND VPWR VPWR U$$1787_1794/HI U$$1787/A1 sky130_fd_sc_hd__conb_1
XFILLER_1_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput220 c[67] VGND VGND VPWR VPWR input220/X sky130_fd_sc_hd__clkbuf_1
Xinput231 c[77] VGND VGND VPWR VPWR input231/X sky130_fd_sc_hd__buf_2
Xinput242 c[87] VGND VGND VPWR VPWR input242/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_3_51_2 dadda_fa_3_51_2/A dadda_fa_3_51_2/B dadda_fa_3_51_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_1/A dadda_fa_4_51_2/B sky130_fd_sc_hd__fa_1
XFILLER_0_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_67_2 U$$939/X U$$1072/X U$$1205/X VGND VGND VPWR VPWR dadda_fa_1_68_6/A
+ dadda_fa_1_67_8/A sky130_fd_sc_hd__fa_1
XFILLER_49_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput253 c[97] VGND VGND VPWR VPWR input253/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_44_1 dadda_fa_3_44_1/A dadda_fa_3_44_1/B dadda_fa_3_44_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_0/CIN dadda_fa_4_44_2/A sky130_fd_sc_hd__fa_1
XFILLER_124_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_21_0 dadda_fa_6_21_0/A dadda_fa_6_21_0/B dadda_fa_6_21_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_22_0/B dadda_fa_7_21_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_37_0 dadda_fa_3_37_0/A dadda_fa_3_37_0/B dadda_fa_3_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_0/B dadda_fa_4_37_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$780 final_adder.U$$780/A final_adder.U$$780/B VGND VGND VPWR VPWR
+ final_adder.U$$780/X sky130_fd_sc_hd__and2_1
XFILLER_75_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$791 final_adder.U$$790/B final_adder.U$$711/X final_adder.U$$679/X
+ VGND VGND VPWR VPWR final_adder.U$$791/X sky130_fd_sc_hd__a21o_1
XU$$630 U$$765/B1 U$$630/A2 U$$632/A1 U$$630/B2 VGND VGND VPWR VPWR U$$631/A sky130_fd_sc_hd__a22o_1
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$641 U$$641/A U$$684/A VGND VGND VPWR VPWR U$$641/X sky130_fd_sc_hd__xor2_1
XFILLER_1_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$652 U$$787/B1 U$$682/A2 U$$654/A1 U$$682/B2 VGND VGND VPWR VPWR U$$653/A sky130_fd_sc_hd__a22o_1
XU$$663 U$$663/A U$$669/B VGND VGND VPWR VPWR U$$663/X sky130_fd_sc_hd__xor2_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$674 U$$811/A1 U$$674/A2 U$$811/B1 U$$674/B2 VGND VGND VPWR VPWR U$$675/A sky130_fd_sc_hd__a22o_1
XU$$685 U$$685/A VGND VGND VPWR VPWR U$$685/Y sky130_fd_sc_hd__inv_1
XU$$696 U$$696/A U$$778/B VGND VGND VPWR VPWR U$$696/X sky130_fd_sc_hd__xor2_1
XFILLER_32_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_96_4 U$$4056/X U$$4189/X U$$4322/X VGND VGND VPWR VPWR dadda_fa_3_97_1/CIN
+ dadda_fa_3_96_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_89_3 input244/X dadda_fa_2_89_3/B dadda_fa_2_89_3/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_90_1/B dadda_fa_3_89_3/B sky130_fd_sc_hd__fa_1
XFILLER_4_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout409 U$$676/A2 VGND VGND VPWR VPWR U$$636/A2 sky130_fd_sc_hd__buf_4
XFILLER_86_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_59_1 dadda_fa_5_59_1/A dadda_fa_5_59_1/B dadda_fa_5_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_60_0/B dadda_fa_7_59_0/A sky130_fd_sc_hd__fa_1
XFILLER_39_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_105_1 U$$3276/X U$$3409/X U$$3542/X VGND VGND VPWR VPWR dadda_fa_3_106_3/B
+ dadda_fa_4_105_0/A sky130_fd_sc_hd__fa_1
XFILLER_81_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2070 U$$2070/A U$$2106/B VGND VGND VPWR VPWR U$$2070/X sky130_fd_sc_hd__xor2_1
XU$$2081 U$$2629/A1 U$$2139/A2 U$$2631/A1 U$$2139/B2 VGND VGND VPWR VPWR U$$2082/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2092 U$$2092/A U$$2096/B VGND VGND VPWR VPWR U$$2092/X sky130_fd_sc_hd__xor2_1
XFILLER_22_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1380 U$$969/A1 U$$1414/A2 U$$3298/B1 U$$1414/B2 VGND VGND VPWR VPWR U$$1381/A
+ sky130_fd_sc_hd__a22o_1
XU$$1391 U$$1391/A U$$1427/B VGND VGND VPWR VPWR U$$1391/X sky130_fd_sc_hd__xor2_1
XFILLER_50_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_84_2 U$$2170/X U$$2303/X U$$2436/X VGND VGND VPWR VPWR dadda_fa_2_85_2/CIN
+ dadda_fa_2_84_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_61_1 dadda_fa_4_61_1/A dadda_fa_4_61_1/B dadda_fa_4_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_62_0/B dadda_fa_5_61_1/B sky130_fd_sc_hd__fa_1
Xfanout910 U$$1202/B2 VGND VGND VPWR VPWR U$$1218/B2 sky130_fd_sc_hd__buf_6
Xfanout921 U$$4508/B2 VGND VGND VPWR VPWR U$$4428/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_77_1 U$$1757/X U$$1890/X U$$2023/X VGND VGND VPWR VPWR dadda_fa_2_78_0/CIN
+ dadda_fa_2_77_3/CIN sky130_fd_sc_hd__fa_1
Xfanout932 fanout938/X VGND VGND VPWR VPWR U$$3376/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_104_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout943 U$$697/B1 VGND VGND VPWR VPWR U$$14/A1 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_4_54_0 dadda_fa_4_54_0/A dadda_fa_4_54_0/B dadda_fa_4_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_55_0/A dadda_fa_5_54_1/A sky130_fd_sc_hd__fa_1
Xfanout954 U$$4470/A1 VGND VGND VPWR VPWR U$$4196/A1 sky130_fd_sc_hd__buf_4
Xfanout965 fanout966/X VGND VGND VPWR VPWR U$$4468/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout976 fanout984/X VGND VGND VPWR VPWR U$$900/B1 sky130_fd_sc_hd__buf_4
XFILLER_86_952 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout987 fanout993/X VGND VGND VPWR VPWR U$$3638/B1 sky130_fd_sc_hd__buf_4
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout998 U$$74/B1 VGND VGND VPWR VPWR U$$76/A1 sky130_fd_sc_hd__buf_4
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_372_ _375_/CLK _372_/D VGND VGND VPWR VPWR _372_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_99_2 dadda_fa_3_99_2/A dadda_fa_3_99_2/B dadda_fa_3_99_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_100_1/A dadda_fa_4_99_2/B sky130_fd_sc_hd__fa_1
XFILLER_126_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_69_0 dadda_fa_6_69_0/A dadda_fa_6_69_0/B dadda_fa_6_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_70_0/B dadda_fa_7_69_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_72_0 dadda_fa_0_72_0/A U$$683/X U$$816/X VGND VGND VPWR VPWR dadda_fa_1_73_7/A
+ dadda_fa_1_72_8/A sky130_fd_sc_hd__fa_1
XFILLER_77_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1006 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$460 U$$460/A U$$498/B VGND VGND VPWR VPWR U$$460/X sky130_fd_sc_hd__xor2_1
XU$$471 U$$882/A1 U$$505/A2 U$$882/B1 U$$505/B2 VGND VGND VPWR VPWR U$$472/A sky130_fd_sc_hd__a22o_1
XU$$482 U$$482/A U$$506/B VGND VGND VPWR VPWR U$$482/X sky130_fd_sc_hd__xor2_1
XU$$493 U$$765/B1 U$$497/A2 U$$632/A1 U$$497/B2 VGND VGND VPWR VPWR U$$494/A sky130_fd_sc_hd__a22o_1
XFILLER_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_94_1 U$$3121/X U$$3254/X U$$3387/X VGND VGND VPWR VPWR dadda_fa_3_95_0/CIN
+ dadda_fa_3_94_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_71_0 dadda_fa_5_71_0/A dadda_fa_5_71_0/B dadda_fa_5_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_72_0/A dadda_fa_6_71_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_87_0 U$$3639/X U$$3772/X U$$3905/X VGND VGND VPWR VPWR dadda_fa_3_88_0/B
+ dadda_fa_3_87_2/B sky130_fd_sc_hd__fa_1
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_70_8 dadda_fa_1_70_8/A dadda_fa_1_70_8/B dadda_fa_1_70_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_71_3/A dadda_fa_3_70_0/A sky130_fd_sc_hd__fa_2
XFILLER_141_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_63_7 dadda_fa_1_63_7/A dadda_fa_1_63_7/B dadda_fa_1_63_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_64_2/CIN dadda_fa_2_63_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_56_6 U$$3577/X U$$3710/X U$$3843/X VGND VGND VPWR VPWR dadda_fa_2_57_2/B
+ dadda_fa_2_56_5/B sky130_fd_sc_hd__fa_1
XFILLER_54_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_49_5 U$$2100/X U$$2233/X U$$2366/X VGND VGND VPWR VPWR dadda_fa_2_50_2/B
+ dadda_fa_2_49_5/B sky130_fd_sc_hd__fa_1
XFILLER_83_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_8_0 dadda_fa_7_8_0/A dadda_fa_7_8_0/B dadda_fa_7_8_0/CIN VGND VGND VPWR
+ VPWR _305_/D _176_/D sky130_fd_sc_hd__fa_1
XFILLER_39_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_86_0 dadda_fa_7_86_0/A dadda_fa_7_86_0/B dadda_fa_7_86_0/CIN VGND VGND
+ VPWR VPWR _383_/D _254_/D sky130_fd_sc_hd__fa_2
XFILLER_109_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1705 fanout1708/X VGND VGND VPWR VPWR U$$4214/B1 sky130_fd_sc_hd__buf_4
XFILLER_105_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1716 U$$4486/B1 VGND VGND VPWR VPWR U$$4488/A1 sky130_fd_sc_hd__buf_2
Xfanout1727 U$$922/A1 VGND VGND VPWR VPWR U$$98/B1 sky130_fd_sc_hd__buf_6
XFILLER_104_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1738 input104/X VGND VGND VPWR VPWR U$$370/B1 sky130_fd_sc_hd__buf_4
Xfanout740 U$$3692/B2 VGND VGND VPWR VPWR U$$3682/B2 sky130_fd_sc_hd__buf_4
Xfanout751 U$$3430/X VGND VGND VPWR VPWR U$$3439/B2 sky130_fd_sc_hd__buf_6
XFILLER_120_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1749 U$$3382/B1 VGND VGND VPWR VPWR U$$4478/B1 sky130_fd_sc_hd__buf_4
Xfanout762 U$$3245/B2 VGND VGND VPWR VPWR U$$3207/B2 sky130_fd_sc_hd__buf_4
XU$$4208 U$$4482/A1 U$$4224/A2 U$$4484/A1 U$$4224/B2 VGND VGND VPWR VPWR U$$4209/A
+ sky130_fd_sc_hd__a22o_1
Xfanout773 U$$3019/X VGND VGND VPWR VPWR U$$3112/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4219 U$$4219/A U$$4231/B VGND VGND VPWR VPWR U$$4219/X sky130_fd_sc_hd__xor2_1
Xfanout784 U$$2882/X VGND VGND VPWR VPWR U$$2989/B2 sky130_fd_sc_hd__buf_2
Xfanout795 U$$279/X VGND VGND VPWR VPWR U$$386/B2 sky130_fd_sc_hd__buf_6
XU$$3507 U$$3642/B1 U$$3511/A2 U$$3509/A1 U$$3511/B2 VGND VGND VPWR VPWR U$$3508/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3518 U$$3518/A U$$3558/B VGND VGND VPWR VPWR U$$3518/X sky130_fd_sc_hd__xor2_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_101_0 dadda_fa_6_101_0/A dadda_fa_6_101_0/B dadda_fa_6_101_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_102_0/B dadda_fa_7_101_0/CIN sky130_fd_sc_hd__fa_1
XU$$3529 U$$4349/B1 U$$3549/A2 U$$4214/B1 U$$3549/B2 VGND VGND VPWR VPWR U$$3530/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2806 U$$4450/A1 U$$2844/A2 U$$4315/A1 U$$2844/B2 VGND VGND VPWR VPWR U$$2807/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2817 U$$2817/A U$$2876/A VGND VGND VPWR VPWR U$$2817/X sky130_fd_sc_hd__xor2_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2828 U$$3239/A1 U$$2840/A2 U$$3239/B1 U$$2840/B2 VGND VGND VPWR VPWR U$$2829/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2839 U$$2839/A U$$2841/B VGND VGND VPWR VPWR U$$2839/X sky130_fd_sc_hd__xor2_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_355_ _356_/CLK _355_/D VGND VGND VPWR VPWR _355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_286_ _421_/CLK _286_/D VGND VGND VPWR VPWR _286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_66_5 dadda_fa_2_66_5/A dadda_fa_2_66_5/B dadda_fa_2_66_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_2/A dadda_fa_4_66_0/A sky130_fd_sc_hd__fa_1
XFILLER_110_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_59_4 dadda_fa_2_59_4/A dadda_fa_2_59_4/B dadda_fa_2_59_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_1/CIN dadda_fa_3_59_3/CIN sky130_fd_sc_hd__fa_1
Xinput6 a[14] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$290 U$$16/A1 U$$312/A2 U$$18/A1 U$$312/B2 VGND VGND VPWR VPWR U$$291/A sky130_fd_sc_hd__a22o_1
XFILLER_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$4 _300_/Q _172_/Q VGND VGND VPWR VPWR final_adder.U$$4/COUT final_adder.U$$4/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_173_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1006 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput310 output310/A VGND VGND VPWR VPWR o[32] sky130_fd_sc_hd__buf_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput321 output321/A VGND VGND VPWR VPWR o[42] sky130_fd_sc_hd__buf_2
Xoutput332 output332/A VGND VGND VPWR VPWR o[52] sky130_fd_sc_hd__buf_2
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 output343/A VGND VGND VPWR VPWR o[62] sky130_fd_sc_hd__buf_2
XFILLER_114_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput354 output354/A VGND VGND VPWR VPWR o[72] sky130_fd_sc_hd__buf_2
Xoutput365 output365/A VGND VGND VPWR VPWR o[82] sky130_fd_sc_hd__buf_2
Xoutput376 output376/A VGND VGND VPWR VPWR o[92] sky130_fd_sc_hd__buf_2
XFILLER_0_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_4 U$$3587/X U$$3720/X U$$3853/X VGND VGND VPWR VPWR dadda_fa_2_62_1/CIN
+ dadda_fa_2_61_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_101_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_3 U$$1977/X U$$2110/X U$$2243/X VGND VGND VPWR VPWR dadda_fa_2_55_1/B
+ dadda_fa_2_54_4/B sky130_fd_sc_hd__fa_1
Xdadda_fa_4_31_2 dadda_fa_4_31_2/A dadda_fa_4_31_2/B dadda_fa_4_31_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_32_0/CIN dadda_fa_5_31_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_47_2 U$$899/X U$$1032/X U$$1165/X VGND VGND VPWR VPWR dadda_fa_2_48_2/A
+ dadda_fa_2_47_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_24_1 dadda_fa_4_24_1/A dadda_fa_4_24_1/B dadda_fa_4_24_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_25_0/B dadda_fa_5_24_1/B sky130_fd_sc_hd__fa_1
XFILLER_83_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_17_0 U$$706/X U$$839/X U$$972/X VGND VGND VPWR VPWR dadda_fa_5_18_0/A
+ dadda_fa_5_17_1/A sky130_fd_sc_hd__fa_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1502 U$$1497/B VGND VGND VPWR VPWR U$$1507/A sky130_fd_sc_hd__buf_6
Xdadda_fa_3_69_3 dadda_fa_3_69_3/A dadda_fa_3_69_3/B dadda_fa_3_69_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_1/B dadda_fa_4_69_2/CIN sky130_fd_sc_hd__fa_1
Xfanout1513 input128/X VGND VGND VPWR VPWR U$$4410/A1 sky130_fd_sc_hd__buf_4
Xfanout1524 U$$981/A1 VGND VGND VPWR VPWR U$$2897/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout1535 U$$979/A1 VGND VGND VPWR VPWR U$$20/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1546 input124/X VGND VGND VPWR VPWR U$$3559/A1 sky130_fd_sc_hd__buf_2
Xfanout1557 U$$4514/A1 VGND VGND VPWR VPWR U$$678/A1 sky130_fd_sc_hd__buf_2
XU$$4005 U$$4416/A1 U$$4005/A2 U$$4416/B1 U$$4005/B2 VGND VGND VPWR VPWR U$$4006/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout570 U$$2272/A2 VGND VGND VPWR VPWR U$$2254/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout1568 input121/X VGND VGND VPWR VPWR U$$4512/A1 sky130_fd_sc_hd__clkbuf_4
XU$$4016 U$$4016/A U$$4098/B VGND VGND VPWR VPWR U$$4016/X sky130_fd_sc_hd__xor2_1
XU$$4027 U$$4162/B1 U$$4045/A2 U$$4027/B1 U$$4045/B2 VGND VGND VPWR VPWR U$$4028/A
+ sky130_fd_sc_hd__a22o_1
Xfanout581 U$$2059/X VGND VGND VPWR VPWR U$$2147/A2 sky130_fd_sc_hd__buf_6
Xfanout1579 U$$3580/A1 VGND VGND VPWR VPWR U$$566/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout592 U$$2022/A2 VGND VGND VPWR VPWR U$$2052/A2 sky130_fd_sc_hd__buf_6
XU$$4038 U$$4038/A U$$4040/B VGND VGND VPWR VPWR U$$4038/X sky130_fd_sc_hd__xor2_1
XU$$4049 U$$4049/A1 U$$4105/A2 U$$4460/B1 U$$4105/B2 VGND VGND VPWR VPWR U$$4050/A
+ sky130_fd_sc_hd__a22o_1
XU$$3304 U$$562/B1 U$$3306/A2 U$$566/A1 U$$3306/B2 VGND VGND VPWR VPWR U$$3305/A sky130_fd_sc_hd__a22o_1
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3315 U$$3315/A U$$3349/B VGND VGND VPWR VPWR U$$3315/X sky130_fd_sc_hd__xor2_1
XU$$3326 U$$4420/B1 U$$3338/A2 U$$4287/A1 U$$3338/B2 VGND VGND VPWR VPWR U$$3327/A
+ sky130_fd_sc_hd__a22o_1
XU$$3337 U$$3337/A U$$3341/B VGND VGND VPWR VPWR U$$3337/X sky130_fd_sc_hd__xor2_1
XFILLER_47_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2603 U$$2603/A VGND VGND VPWR VPWR U$$2603/Y sky130_fd_sc_hd__inv_1
XFILLER_73_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3348 U$$4444/A1 U$$3390/A2 U$$4446/A1 U$$3390/B2 VGND VGND VPWR VPWR U$$3349/A
+ sky130_fd_sc_hd__a22o_1
XU$$3359 U$$3359/A U$$3373/B VGND VGND VPWR VPWR U$$3359/X sky130_fd_sc_hd__xor2_1
XU$$2614 U$$2614/A U$$2668/B VGND VGND VPWR VPWR U$$2614/X sky130_fd_sc_hd__xor2_1
XU$$2625 U$$2625/A1 U$$2665/A2 U$$2762/B1 U$$2665/B2 VGND VGND VPWR VPWR U$$2626/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2636 U$$2636/A U$$2678/B VGND VGND VPWR VPWR U$$2636/X sky130_fd_sc_hd__xor2_1
XU$$1902 U$$1902/A U$$1910/B VGND VGND VPWR VPWR U$$1902/X sky130_fd_sc_hd__xor2_1
XFILLER_92_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2647 U$$2647/A1 U$$2681/A2 U$$183/A1 U$$2681/B2 VGND VGND VPWR VPWR U$$2648/A
+ sky130_fd_sc_hd__a22o_1
XU$$2658 U$$2658/A U$$2662/B VGND VGND VPWR VPWR U$$2658/X sky130_fd_sc_hd__xor2_1
XU$$1913 U$$4377/B1 U$$1915/A2 U$$4244/A1 U$$1915/B2 VGND VGND VPWR VPWR U$$1914/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1924 U$$1924/A1 U$$1964/A2 U$$3022/A1 U$$1964/B2 VGND VGND VPWR VPWR U$$1925/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2669 U$$3628/A1 U$$2711/A2 U$$3628/B1 U$$2711/B2 VGND VGND VPWR VPWR U$$2670/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1935 U$$1935/A U$$1971/B VGND VGND VPWR VPWR U$$1935/X sky130_fd_sc_hd__xor2_1
XU$$1946 U$$2631/A1 U$$1986/A2 U$$2631/B1 U$$1986/B2 VGND VGND VPWR VPWR U$$1947/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1957 U$$1957/A U$$1963/B VGND VGND VPWR VPWR U$$1957/X sky130_fd_sc_hd__xor2_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1968 U$$50/A1 U$$1986/A2 U$$50/B1 U$$1986/B2 VGND VGND VPWR VPWR U$$1969/A sky130_fd_sc_hd__a22o_1
X_407_ _408_/CLK _407_/D VGND VGND VPWR VPWR _407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1979 U$$1979/A U$$2015/B VGND VGND VPWR VPWR U$$1979/X sky130_fd_sc_hd__xor2_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_338_ _338_/CLK _338_/D VGND VGND VPWR VPWR _338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_269_ _408_/CLK _269_/D VGND VGND VPWR VPWR _269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1513_1790 VGND VGND VPWR VPWR U$$1513_1790/HI U$$1513/A1 sky130_fd_sc_hd__conb_1
Xdadda_fa_2_71_3 dadda_fa_2_71_3/A dadda_fa_2_71_3/B dadda_fa_2_71_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_1/B dadda_fa_3_71_3/B sky130_fd_sc_hd__fa_1
Xdadda_fa_2_64_2 dadda_fa_2_64_2/A dadda_fa_2_64_2/B dadda_fa_2_64_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_1/A dadda_fa_3_64_3/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$609 final_adder.U$$608/B final_adder.U$$493/X final_adder.U$$485/X
+ VGND VGND VPWR VPWR final_adder.U$$609/X sky130_fd_sc_hd__a21o_1
XFILLER_97_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_41_1 dadda_fa_5_41_1/A dadda_fa_5_41_1/B dadda_fa_5_41_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_42_0/B dadda_fa_7_41_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_57_1 dadda_fa_2_57_1/A dadda_fa_2_57_1/B dadda_fa_2_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_0/CIN dadda_fa_3_57_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_34_0 dadda_fa_5_34_0/A dadda_fa_5_34_0/B dadda_fa_5_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_35_0/A dadda_fa_6_34_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_110_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$20 U$$20/A1 U$$8/A2 U$$22/A1 U$$8/B2 VGND VGND VPWR VPWR U$$21/A sky130_fd_sc_hd__a22o_1
XU$$31 U$$31/A U$$81/B VGND VGND VPWR VPWR U$$31/X sky130_fd_sc_hd__xor2_1
XU$$42 U$$42/A1 U$$74/A2 U$$44/A1 U$$74/B2 VGND VGND VPWR VPWR U$$43/A sky130_fd_sc_hd__a22o_1
XU$$53 U$$53/A U$$87/B VGND VGND VPWR VPWR U$$53/X sky130_fd_sc_hd__xor2_1
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$64 U$$64/A1 U$$96/A2 U$$64/B1 U$$96/B2 VGND VGND VPWR VPWR U$$65/A sky130_fd_sc_hd__a22o_1
XFILLER_65_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3860 U$$4132/B1 U$$3892/A2 U$$3999/A1 U$$3892/B2 VGND VGND VPWR VPWR U$$3861/A
+ sky130_fd_sc_hd__a22o_1
XU$$75 U$$75/A U$$77/B VGND VGND VPWR VPWR U$$75/X sky130_fd_sc_hd__xor2_1
XU$$3871 U$$3871/A U$$3893/B VGND VGND VPWR VPWR U$$3871/X sky130_fd_sc_hd__xor2_1
XU$$86 U$$86/A1 U$$86/A2 U$$88/A1 U$$86/B2 VGND VGND VPWR VPWR U$$87/A sky130_fd_sc_hd__a22o_1
XU$$3882 U$$4017/B1 U$$3970/A2 U$$3884/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3883/A
+ sky130_fd_sc_hd__a22o_1
XU$$97 U$$97/A U$$97/B VGND VGND VPWR VPWR U$$97/X sky130_fd_sc_hd__xor2_1
XU$$3893 U$$3893/A U$$3893/B VGND VGND VPWR VPWR U$$3893/X sky130_fd_sc_hd__xor2_1
XFILLER_52_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_79_2 dadda_fa_4_79_2/A dadda_fa_4_79_2/B dadda_fa_4_79_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_80_0/CIN dadda_fa_5_79_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_115_971 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_941 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_49_0 dadda_fa_7_49_0/A dadda_fa_7_49_0/B dadda_fa_7_49_0/CIN VGND VGND
+ VPWR VPWR _346_/D _217_/D sky130_fd_sc_hd__fa_1
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_52_0 U$$377/X U$$510/X U$$643/X VGND VGND VPWR VPWR dadda_fa_2_53_0/B
+ dadda_fa_2_52_3/B sky130_fd_sc_hd__fa_1
XFILLER_29_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1209 U$$1209/A U$$1231/B VGND VGND VPWR VPWR U$$1209/X sky130_fd_sc_hd__xor2_1
XFILLER_62_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1003 final_adder.U$$232/A final_adder.U$$733/X final_adder.U$$233/A2
+ VGND VGND VPWR VPWR final_adder.U$$1047/B sky130_fd_sc_hd__a21o_1
XFILLER_8_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1025 final_adder.U$$1/SUM final_adder.U$$255/A2 VGND VGND VPWR VPWR
+ output296/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1036 final_adder.U$$242/A final_adder.U$$623/X VGND VGND VPWR VPWR
+ output288/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1047 final_adder.U$$232/B final_adder.U$$1047/B VGND VGND VPWR VPWR
+ output300/A sky130_fd_sc_hd__xor2_1
XFILLER_109_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1058 final_adder.U$$220/A final_adder.U$$833/X VGND VGND VPWR VPWR
+ output312/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1069 final_adder.U$$210/B final_adder.U$$981/X VGND VGND VPWR VPWR
+ output324/A sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_81_2 dadda_fa_3_81_2/A dadda_fa_3_81_2/B dadda_fa_3_81_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_1/A dadda_fa_4_81_2/B sky130_fd_sc_hd__fa_1
XFILLER_125_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_74_1 dadda_fa_3_74_1/A dadda_fa_3_74_1/B dadda_fa_3_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_0/CIN dadda_fa_4_74_2/A sky130_fd_sc_hd__fa_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_51_0 dadda_fa_6_51_0/A dadda_fa_6_51_0/B dadda_fa_6_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_52_0/B dadda_fa_7_51_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_87_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_67_0 dadda_fa_3_67_0/A dadda_fa_3_67_0/B dadda_fa_3_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_0/B dadda_fa_4_67_1/CIN sky130_fd_sc_hd__fa_1
Xfanout1310 U$$3740/B VGND VGND VPWR VPWR U$$3734/B sky130_fd_sc_hd__buf_6
Xfanout1321 U$$943/B VGND VGND VPWR VPWR U$$959/A sky130_fd_sc_hd__buf_6
XFILLER_87_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1332 U$$3659/B VGND VGND VPWR VPWR U$$3615/B sky130_fd_sc_hd__buf_6
XFILLER_120_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1343 U$$3561/A VGND VGND VPWR VPWR U$$3548/B sky130_fd_sc_hd__buf_6
XFILLER_94_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1354 input44/X VGND VGND VPWR VPWR U$$3391/B sky130_fd_sc_hd__buf_4
Xfanout1365 U$$3073/B VGND VGND VPWR VPWR U$$3061/B sky130_fd_sc_hd__buf_6
Xfanout1376 input38/X VGND VGND VPWR VPWR U$$2974/B sky130_fd_sc_hd__buf_6
XFILLER_4_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1387 U$$2873/B VGND VGND VPWR VPWR U$$2811/B sky130_fd_sc_hd__buf_6
XU$$3101 U$$3101/A U$$3107/B VGND VGND VPWR VPWR U$$3101/X sky130_fd_sc_hd__xor2_1
XFILLER_94_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1398 U$$214/B VGND VGND VPWR VPWR U$$182/B sky130_fd_sc_hd__buf_2
XU$$3112 U$$3112/A1 U$$3112/A2 U$$922/A1 U$$3112/B2 VGND VGND VPWR VPWR U$$3113/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_110_2 dadda_fa_4_110_2/A dadda_fa_4_110_2/B dadda_ha_3_110_3/SUM VGND
+ VGND VPWR VPWR dadda_fa_5_111_0/CIN dadda_fa_5_110_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3123 U$$3123/A U$$3123/B VGND VGND VPWR VPWR U$$3123/X sky130_fd_sc_hd__xor2_1
XU$$3134 U$$3817/B1 U$$3148/A2 U$$3684/A1 U$$3148/B2 VGND VGND VPWR VPWR U$$3135/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2400 U$$2400/A U$$2402/B VGND VGND VPWR VPWR U$$2400/X sky130_fd_sc_hd__xor2_1
XU$$3145 U$$3145/A U$$3147/B VGND VGND VPWR VPWR U$$3145/X sky130_fd_sc_hd__xor2_1
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3156 U$$3154/B U$$3151/A input41/X U$$3151/Y VGND VGND VPWR VPWR U$$3156/X sky130_fd_sc_hd__a22o_2
XU$$2411 U$$82/A1 U$$2415/A2 U$$82/B1 U$$2415/B2 VGND VGND VPWR VPWR U$$2412/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_103_1 dadda_fa_4_103_1/A dadda_fa_4_103_1/B dadda_fa_4_103_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_104_0/B dadda_fa_5_103_1/B sky130_fd_sc_hd__fa_1
XU$$2422 U$$2422/A U$$2456/B VGND VGND VPWR VPWR U$$2422/X sky130_fd_sc_hd__xor2_1
XU$$3167 U$$973/B1 U$$3255/A2 U$$840/A1 U$$3255/B2 VGND VGND VPWR VPWR U$$3168/A sky130_fd_sc_hd__a22o_1
XU$$2433 U$$2707/A1 U$$2443/A2 U$$2707/B1 U$$2443/B2 VGND VGND VPWR VPWR U$$2434/A
+ sky130_fd_sc_hd__a22o_1
XU$$3178 U$$3178/A U$$3210/B VGND VGND VPWR VPWR U$$3178/X sky130_fd_sc_hd__xor2_1
XU$$3189 U$$3189/A1 U$$3199/A2 U$$3189/B1 U$$3199/B2 VGND VGND VPWR VPWR U$$3190/A
+ sky130_fd_sc_hd__a22o_1
XU$$2444 U$$2444/A U$$2446/B VGND VGND VPWR VPWR U$$2444/X sky130_fd_sc_hd__xor2_1
XFILLER_62_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2455 U$$3551/A1 U$$2459/A2 U$$3416/A1 U$$2459/B2 VGND VGND VPWR VPWR U$$2456/A
+ sky130_fd_sc_hd__a22o_1
XU$$1710 U$$749/B1 U$$1720/A2 U$$616/A1 U$$1720/B2 VGND VGND VPWR VPWR U$$1711/A sky130_fd_sc_hd__a22o_1
XU$$2466 U$$2466/A VGND VGND VPWR VPWR U$$2466/Y sky130_fd_sc_hd__inv_1
XU$$1721 U$$1721/A U$$1721/B VGND VGND VPWR VPWR U$$1721/X sky130_fd_sc_hd__xor2_1
XU$$1732 U$$3239/A1 U$$1774/A2 U$$3239/B1 U$$1774/B2 VGND VGND VPWR VPWR U$$1733/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2477 U$$2477/A U$$2545/B VGND VGND VPWR VPWR U$$2477/X sky130_fd_sc_hd__xor2_1
XU$$1504_1789 VGND VGND VPWR VPWR U$$1504_1789/HI U$$1504/B1 sky130_fd_sc_hd__conb_1
XU$$1743 U$$1743/A U$$1761/B VGND VGND VPWR VPWR U$$1743/X sky130_fd_sc_hd__xor2_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2488 U$$2625/A1 U$$2532/A2 U$$2762/B1 U$$2532/B2 VGND VGND VPWR VPWR U$$2489/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2499 U$$2499/A U$$2541/B VGND VGND VPWR VPWR U$$2499/X sky130_fd_sc_hd__xor2_1
XU$$1754 U$$4220/A1 U$$1760/A2 U$$4220/B1 U$$1760/B2 VGND VGND VPWR VPWR U$$1755/A
+ sky130_fd_sc_hd__a22o_1
XU$$1765 U$$1765/A U$$1777/B VGND VGND VPWR VPWR U$$1765/X sky130_fd_sc_hd__xor2_1
XU$$1776 U$$4377/B1 U$$1778/A2 U$$4244/A1 U$$1778/B2 VGND VGND VPWR VPWR U$$1777/A
+ sky130_fd_sc_hd__a22o_1
XU$$1787 U$$1787/A1 U$$1829/A2 U$$3022/A1 U$$1829/B2 VGND VGND VPWR VPWR U$$1788/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1798 U$$1798/A U$$1832/B VGND VGND VPWR VPWR U$$1798/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_124_0 dadda_fa_7_124_0/A dadda_fa_7_124_0/B dadda_fa_7_124_0/CIN VGND
+ VGND VPWR VPWR _421_/D _292_/D sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_41_clk _218_/CLK VGND VGND VPWR VPWR _361_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput20 a[27] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__buf_4
Xinput31 a[37] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput42 a[47] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_1
Xinput53 a[57] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_1
Xinput64 a[9] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_5_89_1 dadda_fa_5_89_1/A dadda_fa_5_89_1/B dadda_fa_5_89_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_90_0/B dadda_fa_7_89_0/A sky130_fd_sc_hd__fa_1
Xinput75 b[19] VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__buf_4
XFILLER_116_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput86 b[29] VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput97 b[39] VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$406 final_adder.U$$410/B final_adder.U$$406/B VGND VGND VPWR VPWR
+ final_adder.U$$530/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$417 final_adder.U$$416/B final_adder.U$$295/X final_adder.U$$291/X
+ VGND VGND VPWR VPWR final_adder.U$$417/X sky130_fd_sc_hd__a21o_1
XFILLER_111_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$428 final_adder.U$$432/B final_adder.U$$428/B VGND VGND VPWR VPWR
+ final_adder.U$$552/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$439 final_adder.U$$438/B final_adder.U$$317/X final_adder.U$$313/X
+ VGND VGND VPWR VPWR final_adder.U$$439/X sky130_fd_sc_hd__a21o_1
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4380 U$$4380/A U$$4383/A VGND VGND VPWR VPWR U$$4380/X sky130_fd_sc_hd__xor2_1
XU$$4391 U$$4391/A U$$4391/B VGND VGND VPWR VPWR U$$4391/X sky130_fd_sc_hd__xor2_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3690 U$$4375/A1 U$$3696/A2 U$$4375/B1 U$$3696/B2 VGND VGND VPWR VPWR U$$3691/A
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_32_clk _388_/CLK VGND VGND VPWR VPWR _386_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_91_1 dadda_fa_4_91_1/A dadda_fa_4_91_1/B dadda_fa_4_91_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_92_0/B dadda_fa_5_91_1/B sky130_fd_sc_hd__fa_1
XFILLER_153_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_84_0 dadda_fa_4_84_0/A dadda_fa_4_84_0/B dadda_fa_4_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_85_0/A dadda_fa_5_84_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_105_3 dadda_fa_3_105_3/A dadda_fa_3_105_3/B dadda_fa_3_105_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_106_1/B dadda_fa_4_105_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$951 final_adder.U$$180/A final_adder.U$$889/X final_adder.U$$951/B1
+ VGND VGND VPWR VPWR final_adder.U$$951/X sky130_fd_sc_hd__a21o_1
XU$$801 U$$936/B1 U$$809/A2 U$$803/A1 U$$809/B2 VGND VGND VPWR VPWR U$$802/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$973 final_adder.U$$202/A final_adder.U$$815/X final_adder.U$$973/B1
+ VGND VGND VPWR VPWR final_adder.U$$973/X sky130_fd_sc_hd__a21o_1
XU$$812 U$$812/A U$$820/B VGND VGND VPWR VPWR U$$812/X sky130_fd_sc_hd__xor2_1
XFILLER_169_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$823 input4/X VGND VGND VPWR VPWR U$$825/B sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$995 final_adder.U$$224/A final_adder.U$$725/X final_adder.U$$995/B1
+ VGND VGND VPWR VPWR final_adder.U$$995/X sky130_fd_sc_hd__a21o_1
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$834 U$$971/A1 U$$904/A2 U$$973/A1 U$$904/B2 VGND VGND VPWR VPWR U$$835/A sky130_fd_sc_hd__a22o_1
XFILLER_28_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$845 U$$845/A U$$875/B VGND VGND VPWR VPWR U$$845/X sky130_fd_sc_hd__xor2_1
XU$$856 U$$856/A1 U$$902/A2 U$$995/A1 U$$902/B2 VGND VGND VPWR VPWR U$$857/A sky130_fd_sc_hd__a22o_1
XU$$867 U$$867/A U$$925/B VGND VGND VPWR VPWR U$$867/X sky130_fd_sc_hd__xor2_1
XU$$1006 U$$1006/A U$$980/B VGND VGND VPWR VPWR U$$1006/X sky130_fd_sc_hd__xor2_1
XU$$1017 U$$56/B1 U$$999/A2 U$$469/B1 U$$999/B2 VGND VGND VPWR VPWR U$$1018/A sky130_fd_sc_hd__a22o_1
XU$$878 U$$878/A1 U$$910/A2 U$$878/B1 U$$910/B2 VGND VGND VPWR VPWR U$$879/A sky130_fd_sc_hd__a22o_1
XFILLER_16_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1028 U$$1028/A U$$998/B VGND VGND VPWR VPWR U$$1028/X sky130_fd_sc_hd__xor2_1
XU$$889 U$$889/A U$$895/B VGND VGND VPWR VPWR U$$889/X sky130_fd_sc_hd__xor2_2
XU$$1039 U$$215/B1 U$$1087/A2 U$$82/A1 U$$1087/B2 VGND VGND VPWR VPWR U$$1040/A sky130_fd_sc_hd__a22o_1
XFILLER_73_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_99_0 dadda_fa_6_99_0/A dadda_fa_6_99_0/B dadda_fa_6_99_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_100_0/B dadda_fa_7_99_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_8_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3979_1828 VGND VGND VPWR VPWR U$$3979_1828/HI U$$3979/A1 sky130_fd_sc_hd__conb_1
XFILLER_112_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1140 U$$3846/A1 VGND VGND VPWR VPWR U$$3435/A1 sky130_fd_sc_hd__buf_2
Xfanout1151 U$$3056/B1 VGND VGND VPWR VPWR U$$866/A1 sky130_fd_sc_hd__buf_4
XFILLER_78_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1162 U$$4424/B1 VGND VGND VPWR VPWR U$$4426/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_94_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1173 U$$40/A1 VGND VGND VPWR VPWR U$$2780/A1 sky130_fd_sc_hd__clkbuf_2
Xfanout1184 input71/X VGND VGND VPWR VPWR U$$4422/A1 sky130_fd_sc_hd__buf_4
Xfanout1195 U$$990/B VGND VGND VPWR VPWR U$$962/A sky130_fd_sc_hd__buf_4
Xdadda_fa_2_41_4 dadda_fa_2_41_4/A dadda_fa_2_41_4/B dadda_fa_2_41_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_42_1/CIN dadda_fa_3_41_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_34_3 U$$1538/X U$$1671/X U$$1804/X VGND VGND VPWR VPWR dadda_fa_3_35_1/B
+ dadda_fa_3_34_3/B sky130_fd_sc_hd__fa_1
XU$$2230 U$$721/B1 U$$2254/A2 U$$999/A1 U$$2254/B2 VGND VGND VPWR VPWR U$$2231/A sky130_fd_sc_hd__a22o_1
XFILLER_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2241 U$$2241/A U$$2249/B VGND VGND VPWR VPWR U$$2241/X sky130_fd_sc_hd__xor2_1
XU$$2252 U$$745/A1 U$$2252/A2 U$$745/B1 U$$2252/B2 VGND VGND VPWR VPWR U$$2253/A sky130_fd_sc_hd__a22o_1
XU$$2263 U$$2263/A U$$2269/B VGND VGND VPWR VPWR U$$2263/X sky130_fd_sc_hd__xor2_1
XU$$2274 U$$3642/B1 U$$2326/A2 U$$3509/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2275/A
+ sky130_fd_sc_hd__a22o_1
XU$$2285 U$$2285/A U$$2327/B VGND VGND VPWR VPWR U$$2285/X sky130_fd_sc_hd__xor2_1
XU$$1540 U$$1540/A U$$1570/B VGND VGND VPWR VPWR U$$1540/X sky130_fd_sc_hd__xor2_1
XU$$2296 U$$2707/A1 U$$2310/A2 U$$2707/B1 U$$2310/B2 VGND VGND VPWR VPWR U$$2297/A
+ sky130_fd_sc_hd__a22o_1
XU$$1551 U$$866/A1 U$$1567/A2 U$$868/A1 U$$1567/B2 VGND VGND VPWR VPWR U$$1552/A sky130_fd_sc_hd__a22o_1
XU$$1562 U$$1562/A U$$1564/B VGND VGND VPWR VPWR U$$1562/X sky130_fd_sc_hd__xor2_1
XFILLER_15_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1573 U$$749/B1 U$$1587/A2 U$$616/A1 U$$1587/B2 VGND VGND VPWR VPWR U$$1574/A sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_14_clk _370_/CLK VGND VGND VPWR VPWR _391_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1584 U$$1584/A U$$1584/B VGND VGND VPWR VPWR U$$1584/X sky130_fd_sc_hd__xor2_1
XU$$1595 U$$499/A1 U$$1641/A2 U$$90/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1596/A sky130_fd_sc_hd__a22o_1
XFILLER_147_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_79_5 U$$3091/X U$$3224/X U$$3357/X VGND VGND VPWR VPWR dadda_fa_2_80_2/A
+ dadda_fa_2_79_5/A sky130_fd_sc_hd__fa_1
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$203 final_adder.U$$202/B final_adder.U$$973/B1 final_adder.U$$203/B1
+ VGND VGND VPWR VPWR final_adder.U$$203/X sky130_fd_sc_hd__a21o_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$214 final_adder.U$$214/A final_adder.U$$214/B VGND VGND VPWR VPWR
+ final_adder.U$$342/B sky130_fd_sc_hd__and2_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$225 final_adder.U$$224/B final_adder.U$$995/B1 final_adder.U$$225/B1
+ VGND VGND VPWR VPWR final_adder.U$$225/X sky130_fd_sc_hd__a21o_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$236 final_adder.U$$236/A final_adder.U$$236/B VGND VGND VPWR VPWR
+ final_adder.U$$364/B sky130_fd_sc_hd__and2_1
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$247 final_adder.U$$9/SUM final_adder.U$$8/COUT final_adder.U$$9/COUT
+ VGND VGND VPWR VPWR final_adder.U$$247/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$258 final_adder.U$$260/B final_adder.U$$258/B VGND VGND VPWR VPWR
+ final_adder.U$$384/B sky130_fd_sc_hd__and2_1
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$269 final_adder.U$$268/B final_adder.U$$143/X final_adder.U$$141/X
+ VGND VGND VPWR VPWR final_adder.U$$269/X sky130_fd_sc_hd__a21o_1
XFILLER_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$108 U$$654/B1 U$$120/A2 U$$521/A1 U$$120/B2 VGND VGND VPWR VPWR U$$109/A sky130_fd_sc_hd__a22o_1
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$119 U$$119/A U$$121/B VGND VGND VPWR VPWR U$$119/X sky130_fd_sc_hd__xor2_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_110_1 U$$3552/X U$$3685/X U$$3818/X VGND VGND VPWR VPWR dadda_fa_4_111_1/A
+ dadda_fa_4_110_2/A sky130_fd_sc_hd__fa_1
XFILLER_119_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_103_0 U$$3937/X U$$4070/X U$$4203/X VGND VGND VPWR VPWR dadda_fa_4_104_0/B
+ dadda_fa_4_103_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_162_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_68_5 U$$2271/X U$$2404/X VGND VGND VPWR VPWR dadda_fa_1_69_7/B dadda_fa_2_68_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput210 c[58] VGND VGND VPWR VPWR input210/X sky130_fd_sc_hd__clkbuf_2
Xinput221 c[68] VGND VGND VPWR VPWR input221/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput232 c[78] VGND VGND VPWR VPWR input232/X sky130_fd_sc_hd__clkbuf_2
Xinput243 c[88] VGND VGND VPWR VPWR input243/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_51_3 dadda_fa_3_51_3/A dadda_fa_3_51_3/B dadda_fa_3_51_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_1/B dadda_fa_4_51_2/CIN sky130_fd_sc_hd__fa_1
Xinput254 c[98] VGND VGND VPWR VPWR input254/X sky130_fd_sc_hd__buf_4
Xdadda_fa_0_67_3 U$$1338/X U$$1471/X U$$1604/X VGND VGND VPWR VPWR dadda_fa_1_68_6/B
+ dadda_fa_1_67_8/B sky130_fd_sc_hd__fa_1
XFILLER_49_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_44_2 dadda_fa_3_44_2/A dadda_fa_3_44_2/B dadda_fa_3_44_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_1/A dadda_fa_4_44_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$770 final_adder.U$$770/A final_adder.U$$770/B VGND VGND VPWR VPWR
+ final_adder.U$$770/X sky130_fd_sc_hd__and2_1
XFILLER_91_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$781 final_adder.U$$780/B final_adder.U$$701/X final_adder.U$$669/X
+ VGND VGND VPWR VPWR final_adder.U$$781/X sky130_fd_sc_hd__a21o_1
XU$$620 U$$70/B1 U$$636/A2 U$$620/B1 U$$636/B2 VGND VGND VPWR VPWR U$$621/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_37_1 dadda_fa_3_37_1/A dadda_fa_3_37_1/B dadda_fa_3_37_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_0/CIN dadda_fa_4_37_2/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$792 final_adder.U$$792/A final_adder.U$$792/B VGND VGND VPWR VPWR
+ final_adder.U$$792/X sky130_fd_sc_hd__and2_1
XU$$631 U$$631/A U$$631/B VGND VGND VPWR VPWR U$$631/X sky130_fd_sc_hd__xor2_1
XFILLER_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$642 U$$916/A1 U$$642/A2 U$$918/A1 U$$642/B2 VGND VGND VPWR VPWR U$$643/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_14_0 dadda_fa_6_14_0/A dadda_fa_6_14_0/B dadda_fa_6_14_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_15_0/B dadda_fa_7_14_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_44_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$653 U$$653/A U$$684/A VGND VGND VPWR VPWR U$$653/X sky130_fd_sc_hd__xor2_1
XU$$664 U$$936/B1 U$$674/A2 U$$803/A1 U$$674/B2 VGND VGND VPWR VPWR U$$665/A sky130_fd_sc_hd__a22o_1
XFILLER_56_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$675 U$$675/A U$$685/A VGND VGND VPWR VPWR U$$675/X sky130_fd_sc_hd__xor2_1
XU$$686 input2/X VGND VGND VPWR VPWR U$$688/B sky130_fd_sc_hd__inv_1
XFILLER_16_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$697 U$$697/A1 U$$743/A2 U$$697/B1 U$$743/B2 VGND VGND VPWR VPWR U$$698/A sky130_fd_sc_hd__a22o_1
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_96_5 U$$4455/X input252/X dadda_fa_2_96_5/CIN VGND VGND VPWR VPWR dadda_fa_3_97_2/A
+ dadda_fa_4_96_0/A sky130_fd_sc_hd__fa_1
XFILLER_126_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_89_4 dadda_fa_2_89_4/A dadda_fa_2_89_4/B dadda_fa_2_89_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_90_1/CIN dadda_fa_3_89_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_3_clk _201_/CLK VGND VGND VPWR VPWR _321_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_32_0 U$$71/X U$$204/X U$$337/X VGND VGND VPWR VPWR dadda_fa_3_33_0/B dadda_fa_3_32_2/B
+ sky130_fd_sc_hd__fa_1
XU$$2060 U$$2058/B U$$2055/A input24/X U$$2055/Y VGND VGND VPWR VPWR U$$2060/X sky130_fd_sc_hd__a22o_4
XFILLER_63_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2071 U$$975/A1 U$$2107/A2 U$$18/A1 U$$2107/B2 VGND VGND VPWR VPWR U$$2072/A sky130_fd_sc_hd__a22o_1
XU$$2082 U$$2082/A U$$2130/B VGND VGND VPWR VPWR U$$2082/X sky130_fd_sc_hd__xor2_1
XU$$2093 U$$997/A1 U$$2097/A2 U$$3189/B1 U$$2097/B2 VGND VGND VPWR VPWR U$$2094/A
+ sky130_fd_sc_hd__a22o_1
XU$$1370 U$$1370/A VGND VGND VPWR VPWR U$$1370/Y sky130_fd_sc_hd__inv_1
XU$$4244_1834 VGND VGND VPWR VPWR U$$4244_1834/HI U$$4244/B1 sky130_fd_sc_hd__conb_1
XU$$1381 U$$1381/A U$$1415/B VGND VGND VPWR VPWR U$$1381/X sky130_fd_sc_hd__xor2_1
XU$$1392 U$$2625/A1 U$$1426/A2 U$$983/A1 U$$1426/B2 VGND VGND VPWR VPWR U$$1393/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_119_0 input150/X dadda_fa_5_119_0/B dadda_fa_5_119_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_6_120_0/A dadda_fa_6_119_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_136_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_84_3 U$$2569/X U$$2702/X U$$2835/X VGND VGND VPWR VPWR dadda_fa_2_85_3/A
+ dadda_fa_2_84_5/A sky130_fd_sc_hd__fa_1
XFILLER_143_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout900 U$$1311/B2 VGND VGND VPWR VPWR U$$1309/B2 sky130_fd_sc_hd__buf_4
XFILLER_132_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout911 U$$1101/X VGND VGND VPWR VPWR U$$1202/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_61_2 dadda_fa_4_61_2/A dadda_fa_4_61_2/B dadda_fa_4_61_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_62_0/CIN dadda_fa_5_61_1/CIN sky130_fd_sc_hd__fa_1
Xfanout922 U$$4508/B2 VGND VGND VPWR VPWR U$$4516/B2 sky130_fd_sc_hd__buf_4
XFILLER_132_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_77_2 U$$2156/X U$$2289/X U$$2422/X VGND VGND VPWR VPWR dadda_fa_2_78_1/A
+ dadda_fa_2_77_4/A sky130_fd_sc_hd__fa_1
Xfanout933 U$$910/A1 VGND VGND VPWR VPWR U$$773/A1 sky130_fd_sc_hd__buf_6
Xfanout944 U$$562/A1 VGND VGND VPWR VPWR U$$697/B1 sky130_fd_sc_hd__buf_2
Xfanout955 U$$908/A1 VGND VGND VPWR VPWR U$$4470/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_4_54_1 dadda_fa_4_54_1/A dadda_fa_4_54_1/B dadda_fa_4_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_55_0/B dadda_fa_5_54_1/B sky130_fd_sc_hd__fa_1
Xfanout966 input96/X VGND VGND VPWR VPWR fanout966/X sky130_fd_sc_hd__buf_8
Xfanout977 fanout984/X VGND VGND VPWR VPWR U$$902/A1 sky130_fd_sc_hd__buf_4
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_31_0 dadda_fa_7_31_0/A dadda_fa_7_31_0/B dadda_fa_7_31_0/CIN VGND VGND
+ VPWR VPWR _328_/D _199_/D sky130_fd_sc_hd__fa_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout988 fanout993/X VGND VGND VPWR VPWR U$$3775/B1 sky130_fd_sc_hd__buf_4
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_47_0 dadda_fa_4_47_0/A dadda_fa_4_47_0/B dadda_fa_4_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_48_0/A dadda_fa_5_47_1/A sky130_fd_sc_hd__fa_1
Xfanout999 fanout999/A VGND VGND VPWR VPWR U$$74/B1 sky130_fd_sc_hd__buf_6
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_371_ _375_/CLK _371_/D VGND VGND VPWR VPWR _371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_99_3 dadda_fa_3_99_3/A dadda_fa_3_99_3/B dadda_fa_3_99_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_100_1/B dadda_fa_4_99_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_170_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1650_1792 VGND VGND VPWR VPWR U$$1650_1792/HI U$$1650/A1 sky130_fd_sc_hd__conb_1
XFILLER_141_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_72_1 U$$949/X U$$1082/X U$$1215/X VGND VGND VPWR VPWR dadda_fa_1_73_7/B
+ dadda_fa_1_72_8/B sky130_fd_sc_hd__fa_1
XFILLER_49_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_65_0 U$$3/A U$$270/X U$$403/X VGND VGND VPWR VPWR dadda_fa_1_66_5/B dadda_fa_1_65_7/B
+ sky130_fd_sc_hd__fa_1
XFILLER_92_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$450 U$$450/A U$$506/B VGND VGND VPWR VPWR U$$450/X sky130_fd_sc_hd__xor2_1
XU$$461 U$$596/B1 U$$497/A2 U$$598/B1 U$$497/B2 VGND VGND VPWR VPWR U$$462/A sky130_fd_sc_hd__a22o_1
XU$$472 U$$472/A U$$506/B VGND VGND VPWR VPWR U$$472/X sky130_fd_sc_hd__xor2_1
XFILLER_45_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$483 U$$894/A1 U$$501/A2 U$$896/A1 U$$501/B2 VGND VGND VPWR VPWR U$$484/A sky130_fd_sc_hd__a22o_1
XU$$494 U$$494/A U$$498/B VGND VGND VPWR VPWR U$$494/X sky130_fd_sc_hd__xor2_1
XFILLER_32_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_94_2 U$$3520/X U$$3653/X U$$3786/X VGND VGND VPWR VPWR dadda_fa_3_95_1/A
+ dadda_fa_3_94_3/A sky130_fd_sc_hd__fa_1
XFILLER_172_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_71_1 dadda_fa_5_71_1/A dadda_fa_5_71_1/B dadda_fa_5_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_72_0/B dadda_fa_7_71_0/A sky130_fd_sc_hd__fa_1
XFILLER_172_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_87_1 U$$4038/X U$$4171/X U$$4304/X VGND VGND VPWR VPWR dadda_fa_3_88_0/CIN
+ dadda_fa_3_87_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_119_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_64_0 dadda_fa_5_64_0/A dadda_fa_5_64_0/B dadda_fa_5_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_65_0/A dadda_fa_6_64_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_141_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_63_8 dadda_fa_1_63_8/A dadda_fa_1_63_8/B dadda_fa_1_63_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_64_3/A dadda_fa_3_63_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_1_56_7 U$$3925/B input208/X dadda_fa_1_56_7/CIN VGND VGND VPWR VPWR dadda_fa_2_57_2/CIN
+ dadda_fa_2_56_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_82_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_49_6 U$$2499/X U$$2632/X U$$2765/X VGND VGND VPWR VPWR dadda_fa_2_50_2/CIN
+ dadda_fa_2_49_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_1_90_3 U$$2980/X U$$3113/X VGND VGND VPWR VPWR dadda_fa_2_91_5/A dadda_fa_3_90_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_149_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_79_0 dadda_fa_7_79_0/A dadda_fa_7_79_0/B dadda_fa_7_79_0/CIN VGND VGND
+ VPWR VPWR _376_/D _247_/D sky130_fd_sc_hd__fa_1
XFILLER_163_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_82_0 dadda_fa_1_82_0/A U$$1368/X U$$1501/X VGND VGND VPWR VPWR dadda_fa_2_83_1/B
+ dadda_fa_2_82_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1706 fanout1708/X VGND VGND VPWR VPWR U$$4490/A1 sky130_fd_sc_hd__buf_2
XFILLER_120_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1717 fanout1718/X VGND VGND VPWR VPWR U$$4486/B1 sky130_fd_sc_hd__buf_6
Xfanout1728 U$$922/A1 VGND VGND VPWR VPWR U$$2840/A1 sky130_fd_sc_hd__buf_4
Xfanout730 U$$3704/X VGND VGND VPWR VPWR U$$3777/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout741 U$$3658/B2 VGND VGND VPWR VPWR U$$3692/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout1739 input104/X VGND VGND VPWR VPWR U$$920/A1 sky130_fd_sc_hd__buf_6
Xfanout752 U$$3293/X VGND VGND VPWR VPWR U$$3338/B2 sky130_fd_sc_hd__buf_4
Xfanout763 U$$3245/B2 VGND VGND VPWR VPWR U$$3241/B2 sky130_fd_sc_hd__buf_4
XFILLER_59_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4209 U$$4209/A U$$4215/B VGND VGND VPWR VPWR U$$4209/X sky130_fd_sc_hd__xor2_1
Xfanout774 U$$3019/X VGND VGND VPWR VPWR U$$3124/B2 sky130_fd_sc_hd__buf_6
Xfanout785 U$$3011/B2 VGND VGND VPWR VPWR U$$3005/B2 sky130_fd_sc_hd__buf_4
Xfanout796 U$$2844/B2 VGND VGND VPWR VPWR U$$2798/B2 sky130_fd_sc_hd__buf_4
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3508 U$$3508/A U$$3562/A VGND VGND VPWR VPWR U$$3508/X sky130_fd_sc_hd__xor2_1
XFILLER_74_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3519 U$$4478/A1 U$$3549/A2 U$$4478/B1 U$$3549/B2 VGND VGND VPWR VPWR U$$3520/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2807 U$$2807/A U$$2877/A VGND VGND VPWR VPWR U$$2807/X sky130_fd_sc_hd__xor2_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2818 U$$4460/B1 U$$2872/A2 U$$3916/A1 U$$2872/B2 VGND VGND VPWR VPWR U$$2819/A
+ sky130_fd_sc_hd__a22o_1
XU$$2829 U$$2829/A U$$2841/B VGND VGND VPWR VPWR U$$2829/X sky130_fd_sc_hd__xor2_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_423_ _423_/CLK _423_/D VGND VGND VPWR VPWR _423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_354_ _356_/CLK _354_/D VGND VGND VPWR VPWR _354_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_285_ _421_/CLK _285_/D VGND VGND VPWR VPWR _285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_81_0 dadda_fa_6_81_0/A dadda_fa_6_81_0/B dadda_fa_6_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_82_0/B dadda_fa_7_81_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_97_0 dadda_fa_3_97_0/A dadda_fa_3_97_0/B dadda_fa_3_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_0/B dadda_fa_4_97_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_59_5 dadda_fa_2_59_5/A dadda_fa_2_59_5/B dadda_fa_2_59_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_2/A dadda_fa_4_59_0/A sky130_fd_sc_hd__fa_2
XFILLER_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 a[15] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_65_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2746_1809 VGND VGND VPWR VPWR U$$2746_1809/HI U$$2746/A1 sky130_fd_sc_hd__conb_1
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$280 U$$280/A1 U$$312/A2 U$$965/B1 U$$312/B2 VGND VGND VPWR VPWR U$$281/A sky130_fd_sc_hd__a22o_1
XFILLER_33_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$291 U$$291/A U$$313/B VGND VGND VPWR VPWR U$$291/X sky130_fd_sc_hd__xor2_1
XFILLER_32_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$5 _301_/Q _173_/Q VGND VGND VPWR VPWR final_adder.U$$5/COUT final_adder.U$$5/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_118_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput300 output300/A VGND VGND VPWR VPWR o[23] sky130_fd_sc_hd__buf_2
Xoutput311 output311/A VGND VGND VPWR VPWR o[33] sky130_fd_sc_hd__buf_2
XFILLER_161_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput322 output322/A VGND VGND VPWR VPWR o[43] sky130_fd_sc_hd__buf_2
Xoutput333 output333/A VGND VGND VPWR VPWR o[53] sky130_fd_sc_hd__buf_2
XFILLER_133_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput344 output344/A VGND VGND VPWR VPWR o[63] sky130_fd_sc_hd__buf_2
XU$$3705_1824 VGND VGND VPWR VPWR U$$3705_1824/HI U$$3705/A1 sky130_fd_sc_hd__conb_1
Xoutput355 output355/A VGND VGND VPWR VPWR o[73] sky130_fd_sc_hd__buf_2
XFILLER_142_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput366 output366/A VGND VGND VPWR VPWR o[83] sky130_fd_sc_hd__buf_2
Xoutput377 output377/A VGND VGND VPWR VPWR o[93] sky130_fd_sc_hd__buf_2
XU$$4471_1883 VGND VGND VPWR VPWR U$$4471_1883/HI U$$4471/B sky130_fd_sc_hd__conb_1
XFILLER_114_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_5 U$$3986/X U$$4119/X input214/X VGND VGND VPWR VPWR dadda_fa_2_62_2/A
+ dadda_fa_2_61_5/A sky130_fd_sc_hd__fa_1
XFILLER_56_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_4 U$$2376/X U$$2509/X U$$2642/X VGND VGND VPWR VPWR dadda_fa_2_55_1/CIN
+ dadda_fa_2_54_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_47_3 U$$1298/X U$$1431/X U$$1564/X VGND VGND VPWR VPWR dadda_fa_2_48_2/B
+ dadda_fa_2_47_5/A sky130_fd_sc_hd__fa_1
XFILLER_71_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_24_2 dadda_fa_4_24_2/A dadda_fa_4_24_2/B dadda_fa_4_24_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_25_0/CIN dadda_fa_5_24_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1024_1917 VGND VGND VPWR VPWR final_adder.U$$1024_1917/HI final_adder.U$$1024/B
+ sky130_fd_sc_hd__conb_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_17_1 U$$1105/X input165/X dadda_fa_4_17_1/CIN VGND VGND VPWR VPWR dadda_fa_5_18_0/B
+ dadda_fa_5_17_1/B sky130_fd_sc_hd__fa_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1503 U$$1475/B VGND VGND VPWR VPWR U$$1497/B sky130_fd_sc_hd__clkbuf_4
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1514 U$$981/B1 VGND VGND VPWR VPWR U$$983/A1 sky130_fd_sc_hd__buf_4
Xfanout1525 U$$981/A1 VGND VGND VPWR VPWR U$$4132/A1 sky130_fd_sc_hd__buf_4
XFILLER_132_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1536 U$$840/B1 VGND VGND VPWR VPWR U$$979/A1 sky130_fd_sc_hd__buf_4
Xfanout1547 U$$4516/A1 VGND VGND VPWR VPWR U$$406/A1 sky130_fd_sc_hd__buf_4
Xfanout560 fanout561/X VGND VGND VPWR VPWR U$$2600/A2 sky130_fd_sc_hd__clkbuf_4
XU$$4006 U$$4006/A U$$4006/B VGND VGND VPWR VPWR U$$4006/X sky130_fd_sc_hd__xor2_1
Xfanout1558 U$$4514/A1 VGND VGND VPWR VPWR U$$4512/B1 sky130_fd_sc_hd__buf_4
Xdadda_ha_3_20_3 U$$1244/X U$$1377/X VGND VGND VPWR VPWR dadda_fa_4_21_1/B dadda_ha_3_20_3/SUM
+ sky130_fd_sc_hd__ha_1
Xfanout571 U$$2196/X VGND VGND VPWR VPWR U$$2272/A2 sky130_fd_sc_hd__buf_6
XFILLER_47_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4017 U$$4152/B1 U$$4105/A2 U$$4017/B1 U$$4105/B2 VGND VGND VPWR VPWR U$$4018/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1569 U$$3964/A1 VGND VGND VPWR VPWR U$$4375/A1 sky130_fd_sc_hd__clkbuf_4
XU$$4028 U$$4028/A U$$4040/B VGND VGND VPWR VPWR U$$4028/X sky130_fd_sc_hd__xor2_1
Xfanout582 U$$2181/A2 VGND VGND VPWR VPWR U$$2177/A2 sky130_fd_sc_hd__buf_6
XU$$4039 U$$4176/A1 U$$4045/A2 U$$4176/B1 U$$4045/B2 VGND VGND VPWR VPWR U$$4040/A
+ sky130_fd_sc_hd__a22o_1
Xfanout593 U$$1922/X VGND VGND VPWR VPWR U$$2022/A2 sky130_fd_sc_hd__buf_4
XFILLER_58_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3305 U$$3305/A U$$3349/B VGND VGND VPWR VPWR U$$3305/X sky130_fd_sc_hd__xor2_1
XFILLER_19_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3316 U$$3999/B1 U$$3340/A2 U$$987/B1 U$$3340/B2 VGND VGND VPWR VPWR U$$3317/A
+ sky130_fd_sc_hd__a22o_1
XU$$3327 U$$3327/A U$$3335/B VGND VGND VPWR VPWR U$$3327/X sky130_fd_sc_hd__xor2_1
XFILLER_46_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3338 U$$3338/A1 U$$3338/A2 U$$735/B1 U$$3338/B2 VGND VGND VPWR VPWR U$$3339/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_100_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2604 input32/X VGND VGND VPWR VPWR U$$2606/B sky130_fd_sc_hd__inv_1
XU$$3349 U$$3349/A U$$3349/B VGND VGND VPWR VPWR U$$3349/X sky130_fd_sc_hd__xor2_1
XU$$2615 U$$3298/B1 U$$2667/A2 U$$4259/B1 U$$2667/B2 VGND VGND VPWR VPWR U$$2616/A
+ sky130_fd_sc_hd__a22o_1
XU$$2626 U$$2626/A U$$2662/B VGND VGND VPWR VPWR U$$2626/X sky130_fd_sc_hd__xor2_1
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2637 U$$32/B1 U$$2679/A2 U$$447/A1 U$$2679/B2 VGND VGND VPWR VPWR U$$2638/A sky130_fd_sc_hd__a22o_1
XU$$1903 U$$2175/B1 U$$1911/A2 U$$2042/A1 U$$1911/B2 VGND VGND VPWR VPWR U$$1904/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2648 U$$2648/A U$$2678/B VGND VGND VPWR VPWR U$$2648/X sky130_fd_sc_hd__xor2_1
XU$$2659 U$$3205/B1 U$$2665/A2 U$$3072/A1 U$$2665/B2 VGND VGND VPWR VPWR U$$2660/A
+ sky130_fd_sc_hd__a22o_1
XU$$1914 U$$1914/A U$$1916/B VGND VGND VPWR VPWR U$$1914/X sky130_fd_sc_hd__xor2_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1925 U$$1925/A U$$1963/B VGND VGND VPWR VPWR U$$1925/X sky130_fd_sc_hd__xor2_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1936 U$$840/A1 U$$1980/A2 U$$840/B1 U$$1980/B2 VGND VGND VPWR VPWR U$$1937/A sky130_fd_sc_hd__a22o_1
XFILLER_15_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1947 U$$1947/A U$$1971/B VGND VGND VPWR VPWR U$$1947/X sky130_fd_sc_hd__xor2_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1958 U$$997/B1 U$$1964/A2 U$$864/A1 U$$1964/B2 VGND VGND VPWR VPWR U$$1959/A sky130_fd_sc_hd__a22o_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_406_ _408_/CLK _406_/D VGND VGND VPWR VPWR _406_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1969 U$$1969/A U$$1971/B VGND VGND VPWR VPWR U$$1969/X sky130_fd_sc_hd__xor2_1
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_337_ _353_/CLK _337_/D VGND VGND VPWR VPWR _337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_268_ _397_/CLK _268_/D VGND VGND VPWR VPWR _268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_199_ _344_/CLK _199_/D VGND VGND VPWR VPWR _199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_71_4 dadda_fa_2_71_4/A dadda_fa_2_71_4/B dadda_fa_2_71_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_1/CIN dadda_fa_3_71_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_64_3 dadda_fa_2_64_3/A dadda_fa_2_64_3/B dadda_fa_2_64_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_1/B dadda_fa_3_64_3/B sky130_fd_sc_hd__fa_1
XFILLER_69_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_57_2 dadda_fa_2_57_2/A dadda_fa_2_57_2/B dadda_fa_2_57_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_1/A dadda_fa_3_57_3/A sky130_fd_sc_hd__fa_2
XFILLER_2_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_34_1 dadda_fa_5_34_1/A dadda_fa_5_34_1/B dadda_fa_5_34_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_35_0/B dadda_fa_7_34_0/A sky130_fd_sc_hd__fa_1
XU$$10 U$$10/A1 U$$8/A2 U$$12/A1 U$$8/B2 VGND VGND VPWR VPWR U$$11/A sky130_fd_sc_hd__a22o_1
XU$$21 U$$21/A U$$9/B VGND VGND VPWR VPWR U$$21/X sky130_fd_sc_hd__xor2_1
XU$$32 U$$32/A1 U$$48/A2 U$$32/B1 U$$48/B2 VGND VGND VPWR VPWR U$$33/A sky130_fd_sc_hd__a22o_1
XFILLER_38_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$43 U$$43/A U$$77/B VGND VGND VPWR VPWR U$$43/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_27_0 dadda_fa_5_27_0/A dadda_fa_5_27_0/B dadda_fa_5_27_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_28_0/A dadda_fa_6_27_0/CIN sky130_fd_sc_hd__fa_1
XU$$3850 U$$4259/B1 U$$3892/A2 U$$3850/B1 U$$3892/B2 VGND VGND VPWR VPWR U$$3851/A
+ sky130_fd_sc_hd__a22o_1
XU$$54 U$$54/A1 U$$86/A2 U$$56/A1 U$$86/B2 VGND VGND VPWR VPWR U$$55/A sky130_fd_sc_hd__a22o_1
XU$$65 U$$65/A U$$97/B VGND VGND VPWR VPWR U$$65/X sky130_fd_sc_hd__xor2_1
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3861 U$$3861/A U$$3867/B VGND VGND VPWR VPWR U$$3861/X sky130_fd_sc_hd__xor2_1
XFILLER_65_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$76 U$$76/A1 U$$80/A2 U$$78/A1 U$$80/B2 VGND VGND VPWR VPWR U$$77/A sky130_fd_sc_hd__a22o_1
XU$$87 U$$87/A U$$87/B VGND VGND VPWR VPWR U$$87/X sky130_fd_sc_hd__xor2_1
XU$$3872 U$$4283/A1 U$$3872/A2 U$$4011/A1 U$$3872/B2 VGND VGND VPWR VPWR U$$3873/A
+ sky130_fd_sc_hd__a22o_1
XU$$3883 U$$3883/A U$$3965/B VGND VGND VPWR VPWR U$$3883/X sky130_fd_sc_hd__xor2_1
XU$$3894 U$$4440/B1 U$$3906/A2 U$$4307/A1 U$$3906/B2 VGND VGND VPWR VPWR U$$3895/A
+ sky130_fd_sc_hd__a22o_1
XU$$98 U$$98/A1 U$$98/A2 U$$98/B1 U$$98/B2 VGND VGND VPWR VPWR U$$99/A sky130_fd_sc_hd__a22o_1
XFILLER_52_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_101_0 dadda_fa_5_101_0/A dadda_fa_5_101_0/B dadda_fa_5_101_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_102_0/A dadda_fa_6_101_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_161_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_983 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_52_1 U$$776/X U$$909/X U$$1042/X VGND VGND VPWR VPWR dadda_fa_2_53_0/CIN
+ dadda_fa_2_52_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_45_0 U$$97/X U$$230/X U$$363/X VGND VGND VPWR VPWR dadda_fa_2_46_2/A dadda_fa_2_45_4/B
+ sky130_fd_sc_hd__fa_1
XFILLER_83_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1015 final_adder.U$$244/A final_adder.U$$625/X final_adder.U$$245/A2
+ VGND VGND VPWR VPWR final_adder.U$$1035/B sky130_fd_sc_hd__a21o_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1026 final_adder.U$$252/A final_adder.U$$255/X VGND VGND VPWR VPWR
+ output307/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1037 final_adder.U$$242/B final_adder.U$$1037/B VGND VGND VPWR VPWR
+ output289/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1048 final_adder.U$$230/A final_adder.U$$731/X VGND VGND VPWR VPWR
+ output301/A sky130_fd_sc_hd__xor2_1
XFILLER_125_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1059 final_adder.U$$220/B final_adder.U$$991/X VGND VGND VPWR VPWR
+ output313/A sky130_fd_sc_hd__xor2_1
XFILLER_152_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_81_3 dadda_fa_3_81_3/A dadda_fa_3_81_3/B dadda_fa_3_81_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_1/B dadda_fa_4_81_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_74_2 dadda_fa_3_74_2/A dadda_fa_3_74_2/B dadda_fa_3_74_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_1/A dadda_fa_4_74_2/B sky130_fd_sc_hd__fa_1
XFILLER_87_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1300 U$$3893/B VGND VGND VPWR VPWR U$$3867/B sky130_fd_sc_hd__buf_6
Xdadda_fa_3_67_1 dadda_fa_3_67_1/A dadda_fa_3_67_1/B dadda_fa_3_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_0/CIN dadda_fa_4_67_2/A sky130_fd_sc_hd__fa_1
Xfanout1311 U$$3740/B VGND VGND VPWR VPWR U$$3774/B sky130_fd_sc_hd__buf_6
Xfanout1322 U$$955/B VGND VGND VPWR VPWR U$$943/B sky130_fd_sc_hd__buf_4
Xfanout1333 U$$3698/A VGND VGND VPWR VPWR U$$3695/B sky130_fd_sc_hd__buf_6
Xdadda_fa_6_44_0 dadda_fa_6_44_0/A dadda_fa_6_44_0/B dadda_fa_6_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_45_0/B dadda_fa_7_44_0/CIN sky130_fd_sc_hd__fa_1
Xfanout1344 U$$3524/B VGND VGND VPWR VPWR U$$3561/A sky130_fd_sc_hd__buf_4
Xfanout1355 U$$3208/B VGND VGND VPWR VPWR U$$3196/B sky130_fd_sc_hd__buf_6
Xfanout1366 input40/X VGND VGND VPWR VPWR U$$3073/B sky130_fd_sc_hd__buf_6
Xfanout1377 input38/X VGND VGND VPWR VPWR U$$3014/A sky130_fd_sc_hd__buf_4
Xfanout1388 U$$2876/A VGND VGND VPWR VPWR U$$2871/B sky130_fd_sc_hd__buf_6
XFILLER_59_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout390 U$$1087/A2 VGND VGND VPWR VPWR U$$1093/A2 sky130_fd_sc_hd__buf_6
XU$$3102 U$$3239/A1 U$$3108/A2 U$$3239/B1 U$$3108/B2 VGND VGND VPWR VPWR U$$3103/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1399 U$$210/B VGND VGND VPWR VPWR U$$214/B sky130_fd_sc_hd__clkbuf_4
XU$$3113 U$$3113/A U$$3151/A VGND VGND VPWR VPWR U$$3113/X sky130_fd_sc_hd__xor2_1
XU$$3124 U$$384/A1 U$$3124/A2 U$$384/B1 U$$3124/B2 VGND VGND VPWR VPWR U$$3125/A sky130_fd_sc_hd__a22o_1
XU$$3135 U$$3135/A U$$3150/A VGND VGND VPWR VPWR U$$3135/X sky130_fd_sc_hd__xor2_1
XU$$2401 U$$70/B1 U$$2445/A2 U$$620/B1 U$$2445/B2 VGND VGND VPWR VPWR U$$2402/A sky130_fd_sc_hd__a22o_1
XU$$3146 U$$3418/B1 U$$3148/A2 U$$3285/A1 U$$3148/B2 VGND VGND VPWR VPWR U$$3147/A
+ sky130_fd_sc_hd__a22o_1
XU$$3157 U$$3157/A1 U$$3199/A2 U$$4392/A1 U$$3199/B2 VGND VGND VPWR VPWR U$$3158/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2412 U$$2412/A U$$2412/B VGND VGND VPWR VPWR U$$2412/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_103_2 dadda_fa_4_103_2/A dadda_fa_4_103_2/B dadda_fa_4_103_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_104_0/CIN dadda_fa_5_103_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_34_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2423 U$$3382/A1 U$$2459/A2 U$$3382/B1 U$$2459/B2 VGND VGND VPWR VPWR U$$2424/A
+ sky130_fd_sc_hd__a22o_1
XU$$3168 U$$3168/A U$$3210/B VGND VGND VPWR VPWR U$$3168/X sky130_fd_sc_hd__xor2_1
XU$$2434 U$$2434/A U$$2466/A VGND VGND VPWR VPWR U$$2434/X sky130_fd_sc_hd__xor2_1
XU$$3179 U$$4412/A1 U$$3255/A2 U$$4414/A1 U$$3255/B2 VGND VGND VPWR VPWR U$$3180/A
+ sky130_fd_sc_hd__a22o_1
XU$$1700 U$$56/A1 U$$1702/A2 U$$56/B1 U$$1702/B2 VGND VGND VPWR VPWR U$$1701/A sky130_fd_sc_hd__a22o_1
XU$$2445 U$$938/A1 U$$2445/A2 U$$940/A1 U$$2445/B2 VGND VGND VPWR VPWR U$$2446/A sky130_fd_sc_hd__a22o_1
XU$$1711 U$$1711/A U$$1721/B VGND VGND VPWR VPWR U$$1711/X sky130_fd_sc_hd__xor2_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2456 U$$2456/A U$$2456/B VGND VGND VPWR VPWR U$$2456/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2467 input30/X VGND VGND VPWR VPWR U$$2469/B sky130_fd_sc_hd__inv_1
XU$$1722 U$$900/A1 U$$1726/A2 U$$900/B1 U$$1726/B2 VGND VGND VPWR VPWR U$$1723/A sky130_fd_sc_hd__a22o_1
XU$$4381_1836 VGND VGND VPWR VPWR U$$4381_1836/HI U$$4381/B1 sky130_fd_sc_hd__conb_1
XU$$1733 U$$1733/A U$$1741/B VGND VGND VPWR VPWR U$$1733/X sky130_fd_sc_hd__xor2_1
XU$$2478 U$$3298/B1 U$$2546/A2 U$$2480/A1 U$$2546/B2 VGND VGND VPWR VPWR U$$2479/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2489 U$$2489/A U$$2529/B VGND VGND VPWR VPWR U$$2489/X sky130_fd_sc_hd__xor2_1
XU$$1744 U$$920/B1 U$$1758/A2 U$$787/A1 U$$1758/B2 VGND VGND VPWR VPWR U$$1745/A sky130_fd_sc_hd__a22o_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1755 U$$1755/A U$$1761/B VGND VGND VPWR VPWR U$$1755/X sky130_fd_sc_hd__xor2_1
XU$$1766 U$$2175/B1 U$$1778/A2 U$$2042/A1 U$$1778/B2 VGND VGND VPWR VPWR U$$1767/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1777 U$$1777/A U$$1777/B VGND VGND VPWR VPWR U$$1777/X sky130_fd_sc_hd__xor2_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1788 U$$1788/A U$$1828/B VGND VGND VPWR VPWR U$$1788/X sky130_fd_sc_hd__xor2_1
XFILLER_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1799 U$$3030/B1 U$$1841/A2 U$$2897/A1 U$$1841/B2 VGND VGND VPWR VPWR U$$1800/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_117_0 dadda_fa_7_117_0/A dadda_fa_7_117_0/B dadda_fa_7_117_0/CIN VGND
+ VGND VPWR VPWR _414_/D _285_/D sky130_fd_sc_hd__fa_1
XFILLER_174_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput10 a[18] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_2
Xinput21 a[28] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_1
Xinput32 a[38] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 a[48] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput54 a[58] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_1
Xinput65 b[0] VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__clkbuf_4
Xinput76 b[1] VGND VGND VPWR VPWR input76/X sky130_fd_sc_hd__buf_4
Xinput87 b[2] VGND VGND VPWR VPWR input87/X sky130_fd_sc_hd__clkbuf_2
Xinput98 b[3] VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_62_0 dadda_fa_2_62_0/A dadda_fa_2_62_0/B dadda_fa_2_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_0/B dadda_fa_3_62_2/B sky130_fd_sc_hd__fa_1
XFILLER_96_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$407 final_adder.U$$406/B final_adder.U$$285/X final_adder.U$$281/X
+ VGND VGND VPWR VPWR final_adder.U$$407/X sky130_fd_sc_hd__a21o_1
XFILLER_112_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$418 final_adder.U$$422/B final_adder.U$$418/B VGND VGND VPWR VPWR
+ final_adder.U$$542/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$429 final_adder.U$$428/B final_adder.U$$307/X final_adder.U$$303/X
+ VGND VGND VPWR VPWR final_adder.U$$429/X sky130_fd_sc_hd__a21o_1
XFILLER_84_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4370 U$$4370/A U$$4374/B VGND VGND VPWR VPWR U$$4370/X sky130_fd_sc_hd__xor2_1
XU$$4381 U$$545/A1 U$$4381/A2 U$$4381/B1 U$$4381/B2 VGND VGND VPWR VPWR U$$4382/A
+ sky130_fd_sc_hd__a22o_1
XU$$4392 U$$4392/A1 U$$4388/X input76/X U$$4428/B2 VGND VGND VPWR VPWR U$$4393/A sky130_fd_sc_hd__a22o_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3680 U$$3817/A1 U$$3682/A2 U$$3817/B1 U$$3682/B2 VGND VGND VPWR VPWR U$$3681/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3691 U$$3691/A U$$3695/B VGND VGND VPWR VPWR U$$3691/X sky130_fd_sc_hd__xor2_1
XFILLER_80_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2990 U$$2990/A U$$2990/B VGND VGND VPWR VPWR U$$2990/X sky130_fd_sc_hd__xor2_1
XFILLER_52_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_91_2 dadda_fa_4_91_2/A dadda_fa_4_91_2/B dadda_fa_4_91_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_92_0/CIN dadda_fa_5_91_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_84_1 dadda_fa_4_84_1/A dadda_fa_4_84_1/B dadda_fa_4_84_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_85_0/B dadda_fa_5_84_1/B sky130_fd_sc_hd__fa_1
XFILLER_134_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_61_0 dadda_fa_7_61_0/A dadda_fa_7_61_0/B dadda_fa_7_61_0/CIN VGND VGND
+ VPWR VPWR _358_/D _229_/D sky130_fd_sc_hd__fa_1
XFILLER_162_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_77_0 dadda_fa_4_77_0/A dadda_fa_4_77_0/B dadda_fa_4_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_78_0/A dadda_fa_5_77_1/A sky130_fd_sc_hd__fa_1
XFILLER_106_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_920 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$941 final_adder.U$$170/A final_adder.U$$879/X final_adder.U$$941/B1
+ VGND VGND VPWR VPWR final_adder.U$$941/X sky130_fd_sc_hd__a21o_1
XFILLER_29_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$963 final_adder.U$$192/A final_adder.U$$805/X final_adder.U$$963/B1
+ VGND VGND VPWR VPWR final_adder.U$$963/X sky130_fd_sc_hd__a21o_1
XFILLER_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$802 U$$802/A U$$804/B VGND VGND VPWR VPWR U$$802/X sky130_fd_sc_hd__xor2_1
XU$$813 U$$950/A1 U$$817/A2 U$$952/A1 U$$817/B2 VGND VGND VPWR VPWR U$$814/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$985 final_adder.U$$214/A final_adder.U$$827/X final_adder.U$$985/B1
+ VGND VGND VPWR VPWR final_adder.U$$985/X sky130_fd_sc_hd__a21o_1
XU$$824 U$$959/A VGND VGND VPWR VPWR U$$824/Y sky130_fd_sc_hd__inv_1
XFILLER_84_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$835 U$$835/A U$$907/B VGND VGND VPWR VPWR U$$835/X sky130_fd_sc_hd__xor2_1
XFILLER_90_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$846 U$$24/A1 U$$876/A2 U$$26/A1 U$$876/B2 VGND VGND VPWR VPWR U$$847/A sky130_fd_sc_hd__a22o_1
XU$$857 U$$857/A U$$895/B VGND VGND VPWR VPWR U$$857/X sky130_fd_sc_hd__xor2_1
XFILLER_28_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$868 U$$868/A1 U$$902/A2 U$$868/B1 U$$902/B2 VGND VGND VPWR VPWR U$$869/A sky130_fd_sc_hd__a22o_1
XFILLER_113_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1007 U$$48/A1 U$$979/A2 U$$50/A1 U$$979/B2 VGND VGND VPWR VPWR U$$1008/A sky130_fd_sc_hd__a22o_1
XU$$1018 U$$1018/A U$$1062/B VGND VGND VPWR VPWR U$$1018/X sky130_fd_sc_hd__xor2_1
XU$$879 U$$879/A U$$913/B VGND VGND VPWR VPWR U$$879/X sky130_fd_sc_hd__xor2_1
XU$$1029 U$$892/A1 U$$999/A2 U$$894/A1 U$$999/B2 VGND VGND VPWR VPWR U$$1030/A sky130_fd_sc_hd__a22o_1
XFILLER_19_1042 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1130 U$$3884/A1 VGND VGND VPWR VPWR U$$870/A1 sky130_fd_sc_hd__buf_4
Xfanout1141 input76/X VGND VGND VPWR VPWR U$$3846/A1 sky130_fd_sc_hd__buf_4
XFILLER_152_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1152 U$$4291/A1 VGND VGND VPWR VPWR U$$3056/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1163 U$$40/B1 VGND VGND VPWR VPWR U$$42/A1 sky130_fd_sc_hd__buf_4
XFILLER_94_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1174 U$$4150/A1 VGND VGND VPWR VPWR U$$40/A1 sky130_fd_sc_hd__buf_4
Xfanout1185 U$$3322/B1 VGND VGND VPWR VPWR U$$995/A1 sky130_fd_sc_hd__buf_4
Xfanout1196 input7/X VGND VGND VPWR VPWR U$$990/B sky130_fd_sc_hd__buf_8
Xdadda_fa_2_41_5 dadda_fa_2_41_5/A dadda_fa_2_41_5/B dadda_fa_2_41_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_42_2/A dadda_fa_4_41_0/A sky130_fd_sc_hd__fa_1
XFILLER_47_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2220 U$$850/A1 U$$2254/A2 U$$989/A1 U$$2254/B2 VGND VGND VPWR VPWR U$$2221/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_34_4 U$$1937/X U$$2070/X U$$2203/X VGND VGND VPWR VPWR dadda_fa_3_35_1/CIN
+ dadda_fa_3_34_3/CIN sky130_fd_sc_hd__fa_1
XU$$2231 U$$2231/A U$$2231/B VGND VGND VPWR VPWR U$$2231/X sky130_fd_sc_hd__xor2_1
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2242 U$$872/A1 U$$2248/A2 U$$874/A1 U$$2248/B2 VGND VGND VPWR VPWR U$$2243/A sky130_fd_sc_hd__a22o_1
XU$$2253 U$$2253/A U$$2253/B VGND VGND VPWR VPWR U$$2253/X sky130_fd_sc_hd__xor2_1
XU$$2264 U$$3495/B1 U$$2196/X U$$3499/A1 U$$2197/X VGND VGND VPWR VPWR U$$2265/A sky130_fd_sc_hd__a22o_1
XU$$1530 U$$1530/A U$$1568/B VGND VGND VPWR VPWR U$$1530/X sky130_fd_sc_hd__xor2_1
XU$$2275 U$$2275/A U$$2327/B VGND VGND VPWR VPWR U$$2275/X sky130_fd_sc_hd__xor2_1
XFILLER_16_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1541 U$$32/B1 U$$1587/A2 U$$447/A1 U$$1587/B2 VGND VGND VPWR VPWR U$$1542/A sky130_fd_sc_hd__a22o_1
XU$$2286 U$$4478/A1 U$$2326/A2 U$$4478/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2287/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2297 U$$2297/A U$$2301/B VGND VGND VPWR VPWR U$$2297/X sky130_fd_sc_hd__xor2_1
XU$$1552 U$$1552/A U$$1568/B VGND VGND VPWR VPWR U$$1552/X sky130_fd_sc_hd__xor2_1
XU$$1563 U$$56/A1 U$$1563/A2 U$$56/B1 U$$1563/B2 VGND VGND VPWR VPWR U$$1564/A sky130_fd_sc_hd__a22o_1
XU$$1574 U$$1574/A U$$1584/B VGND VGND VPWR VPWR U$$1574/X sky130_fd_sc_hd__xor2_1
XU$$1585 U$$215/A1 U$$1587/A2 U$$215/B1 U$$1587/B2 VGND VGND VPWR VPWR U$$1586/A sky130_fd_sc_hd__a22o_1
XU$$1596 U$$1596/A U$$1608/B VGND VGND VPWR VPWR U$$1596/X sky130_fd_sc_hd__xor2_1
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_94_0 dadda_fa_5_94_0/A dadda_fa_5_94_0/B dadda_fa_5_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_95_0/A dadda_fa_6_94_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_79_6 U$$3490/X U$$3623/X U$$3756/X VGND VGND VPWR VPWR dadda_fa_2_80_2/B
+ dadda_fa_2_79_5/B sky130_fd_sc_hd__fa_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$204 final_adder.U$$204/A final_adder.U$$204/B VGND VGND VPWR VPWR
+ final_adder.U$$332/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$215 final_adder.U$$214/B final_adder.U$$985/B1 final_adder.U$$215/B1
+ VGND VGND VPWR VPWR final_adder.U$$215/X sky130_fd_sc_hd__a21o_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$226 final_adder.U$$226/A final_adder.U$$226/B VGND VGND VPWR VPWR
+ final_adder.U$$354/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$237 final_adder.U$$236/B final_adder.U$$237/A2 final_adder.U$$237/B1
+ VGND VGND VPWR VPWR final_adder.U$$237/X sky130_fd_sc_hd__a21o_1
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$248 final_adder.U$$6/SUM final_adder.U$$7/SUM VGND VGND VPWR VPWR
+ final_adder.U$$376/B sky130_fd_sc_hd__and2_1
XFILLER_85_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$259 final_adder.U$$258/B final_adder.U$$133/X final_adder.U$$131/X
+ VGND VGND VPWR VPWR final_adder.U$$259/X sky130_fd_sc_hd__a21o_1
XU$$109 U$$109/A U$$121/B VGND VGND VPWR VPWR U$$109/X sky130_fd_sc_hd__xor2_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_951 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4405_1850 VGND VGND VPWR VPWR U$$4405_1850/HI U$$4405/B sky130_fd_sc_hd__conb_1
XFILLER_166_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_110_2 U$$3951/X U$$4084/X U$$4217/X VGND VGND VPWR VPWR dadda_fa_4_111_1/B
+ dadda_fa_4_110_2/B sky130_fd_sc_hd__fa_1
XFILLER_104_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_103_1 U$$4336/X U$$4469/X input133/X VGND VGND VPWR VPWR dadda_fa_4_104_0/CIN
+ dadda_fa_4_103_2/A sky130_fd_sc_hd__fa_1
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput200 c[49] VGND VGND VPWR VPWR input200/X sky130_fd_sc_hd__clkbuf_2
Xinput211 c[59] VGND VGND VPWR VPWR input211/X sky130_fd_sc_hd__clkbuf_2
Xinput222 c[69] VGND VGND VPWR VPWR input222/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_124_0 dadda_fa_6_124_0/A dadda_fa_6_124_0/B dadda_fa_6_124_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_125_0/B dadda_fa_7_124_0/CIN sky130_fd_sc_hd__fa_1
Xinput233 c[79] VGND VGND VPWR VPWR input233/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput244 c[89] VGND VGND VPWR VPWR input244/X sky130_fd_sc_hd__buf_2
Xinput255 c[99] VGND VGND VPWR VPWR input255/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_0_67_4 U$$1737/X U$$1870/X U$$2003/X VGND VGND VPWR VPWR dadda_fa_1_68_6/CIN
+ dadda_fa_1_67_8/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_44_3 dadda_fa_3_44_3/A dadda_fa_3_44_3/B dadda_fa_3_44_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_1/B dadda_fa_4_44_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$760 final_adder.U$$792/B final_adder.U$$760/B VGND VGND VPWR VPWR
+ final_adder.U$$760/X sky130_fd_sc_hd__and2_1
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$771 final_adder.U$$770/B final_adder.U$$691/X final_adder.U$$659/X
+ VGND VGND VPWR VPWR final_adder.U$$771/X sky130_fd_sc_hd__a21o_1
XFILLER_90_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$610 U$$745/B1 U$$610/A2 U$$747/B1 U$$610/B2 VGND VGND VPWR VPWR U$$611/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$782 final_adder.U$$782/A final_adder.U$$782/B VGND VGND VPWR VPWR
+ final_adder.U$$782/X sky130_fd_sc_hd__and2_1
XU$$621 U$$621/A U$$637/B VGND VGND VPWR VPWR U$$621/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_37_2 dadda_fa_3_37_2/A dadda_fa_3_37_2/B dadda_fa_3_37_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_1/A dadda_fa_4_37_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$793 final_adder.U$$792/B final_adder.U$$713/X final_adder.U$$681/X
+ VGND VGND VPWR VPWR final_adder.U$$793/X sky130_fd_sc_hd__a21o_1
XU$$632 U$$632/A1 U$$674/A2 U$$632/B1 U$$674/B2 VGND VGND VPWR VPWR U$$633/A sky130_fd_sc_hd__a22o_1
XFILLER_17_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$643 U$$643/A U$$643/B VGND VGND VPWR VPWR U$$643/X sky130_fd_sc_hd__xor2_1
XU$$654 U$$654/A1 U$$682/A2 U$$654/B1 U$$682/B2 VGND VGND VPWR VPWR U$$655/A sky130_fd_sc_hd__a22o_1
XFILLER_17_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$665 U$$665/A U$$669/B VGND VGND VPWR VPWR U$$665/X sky130_fd_sc_hd__xor2_1
XFILLER_56_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$676 U$$811/B1 U$$676/A2 U$$678/A1 U$$676/B2 VGND VGND VPWR VPWR U$$677/A sky130_fd_sc_hd__a22o_1
XU$$687 U$$804/B VGND VGND VPWR VPWR U$$687/Y sky130_fd_sc_hd__inv_1
XFILLER_17_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$698 U$$698/A U$$744/B VGND VGND VPWR VPWR U$$698/X sky130_fd_sc_hd__xor2_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3842_1826 VGND VGND VPWR VPWR U$$3842_1826/HI U$$3842/A1 sky130_fd_sc_hd__conb_1
XFILLER_144_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_89_5 dadda_fa_2_89_5/A dadda_fa_2_89_5/B dadda_fa_2_89_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_90_2/A dadda_fa_4_89_0/A sky130_fd_sc_hd__fa_1
XFILLER_141_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_2_26_2 U$$857/X U$$990/X VGND VGND VPWR VPWR dadda_fa_3_27_3/A dadda_fa_4_26_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_67_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_32_1 U$$470/X U$$603/X U$$736/X VGND VGND VPWR VPWR dadda_fa_3_33_0/CIN
+ dadda_fa_3_32_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_25_0 U$$57/X U$$190/X U$$323/X VGND VGND VPWR VPWR dadda_fa_3_26_2/CIN
+ dadda_fa_3_25_3/CIN sky130_fd_sc_hd__fa_1
XU$$2050 U$$4377/B1 U$$2052/A2 U$$4244/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2051/A
+ sky130_fd_sc_hd__a22o_1
XU$$2061 U$$2061/A1 U$$2097/A2 U$$3022/A1 U$$2097/B2 VGND VGND VPWR VPWR U$$2062/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2072 U$$2072/A U$$2106/B VGND VGND VPWR VPWR U$$2072/X sky130_fd_sc_hd__xor2_1
XFILLER_23_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2083 U$$2631/A1 U$$2097/A2 U$$2631/B1 U$$2097/B2 VGND VGND VPWR VPWR U$$2084/A
+ sky130_fd_sc_hd__a22o_1
XU$$2094 U$$2094/A U$$2096/B VGND VGND VPWR VPWR U$$2094/X sky130_fd_sc_hd__xor2_1
XU$$1360 U$$1360/A U$$1360/B VGND VGND VPWR VPWR U$$1360/X sky130_fd_sc_hd__xor2_1
XU$$1371 input13/X VGND VGND VPWR VPWR U$$1373/B sky130_fd_sc_hd__inv_1
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1382 U$$3298/B1 U$$1414/A2 U$$2480/A1 U$$1414/B2 VGND VGND VPWR VPWR U$$1383/A
+ sky130_fd_sc_hd__a22o_1
XU$$1393 U$$1393/A U$$1427/B VGND VGND VPWR VPWR U$$1393/X sky130_fd_sc_hd__xor2_1
XFILLER_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_119_1 dadda_fa_5_119_1/A dadda_fa_5_119_1/B dadda_fa_5_119_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_120_0/B dadda_fa_7_119_0/A sky130_fd_sc_hd__fa_1
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4435_1865 VGND VGND VPWR VPWR U$$4435_1865/HI U$$4435/B sky130_fd_sc_hd__conb_1
Xdadda_fa_1_84_4 U$$2968/X U$$3101/X U$$3234/X VGND VGND VPWR VPWR dadda_fa_2_85_3/B
+ dadda_fa_2_84_5/B sky130_fd_sc_hd__fa_1
XFILLER_1_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout901 U$$1353/B2 VGND VGND VPWR VPWR U$$1311/B2 sky130_fd_sc_hd__buf_4
Xfanout912 U$$102/B2 VGND VGND VPWR VPWR U$$96/B2 sky130_fd_sc_hd__buf_4
Xfanout923 U$$4389/X VGND VGND VPWR VPWR U$$4508/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_131_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_77_3 U$$2555/X U$$2688/X U$$2821/X VGND VGND VPWR VPWR dadda_fa_2_78_1/B
+ dadda_fa_2_77_4/B sky130_fd_sc_hd__fa_1
Xfanout934 U$$3650/A1 VGND VGND VPWR VPWR U$$4196/B1 sky130_fd_sc_hd__buf_4
Xfanout945 U$$973/A1 VGND VGND VPWR VPWR U$$562/A1 sky130_fd_sc_hd__buf_2
XFILLER_98_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout956 fanout957/X VGND VGND VPWR VPWR U$$908/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_54_2 dadda_fa_4_54_2/A dadda_fa_4_54_2/B dadda_fa_4_54_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_55_0/CIN dadda_fa_5_54_1/CIN sky130_fd_sc_hd__fa_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout967 fanout975/X VGND VGND VPWR VPWR U$$765/B1 sky130_fd_sc_hd__buf_4
XFILLER_100_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout978 U$$3642/A1 VGND VGND VPWR VPWR U$$3503/B1 sky130_fd_sc_hd__buf_4
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout989 U$$215/A1 VGND VGND VPWR VPWR U$$78/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_47_1 dadda_fa_4_47_1/A dadda_fa_4_47_1/B dadda_fa_4_47_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_48_0/B dadda_fa_5_47_1/B sky130_fd_sc_hd__fa_1
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_24_0 dadda_fa_7_24_0/A dadda_fa_7_24_0/B dadda_fa_7_24_0/CIN VGND VGND
+ VPWR VPWR _321_/D _192_/D sky130_fd_sc_hd__fa_2
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_370_ _370_/CLK _370_/D VGND VGND VPWR VPWR _370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_114_0_1938 VGND VGND VPWR VPWR dadda_fa_3_114_0/A dadda_fa_3_114_0_1938/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_72_2 U$$1348/X U$$1481/X U$$1614/X VGND VGND VPWR VPWR dadda_fa_1_73_7/CIN
+ dadda_fa_1_72_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_65_1 U$$536/X U$$669/X U$$802/X VGND VGND VPWR VPWR dadda_fa_1_66_5/CIN
+ dadda_fa_1_65_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_92_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_42_0 dadda_fa_3_42_0/A dadda_fa_3_42_0/B dadda_fa_3_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_0/B dadda_fa_4_42_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_58_0 U$$123/X U$$256/X U$$389/X VGND VGND VPWR VPWR dadda_fa_1_59_6/CIN
+ dadda_fa_1_58_8/A sky130_fd_sc_hd__fa_1
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$590 final_adder.U$$598/B final_adder.U$$590/B VGND VGND VPWR VPWR
+ final_adder.U$$710/B sky130_fd_sc_hd__and2_1
XFILLER_17_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$440 U$$440/A U$$506/B VGND VGND VPWR VPWR U$$440/X sky130_fd_sc_hd__xor2_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$451 U$$999/A1 U$$501/A2 U$$999/B1 U$$501/B2 VGND VGND VPWR VPWR U$$452/A sky130_fd_sc_hd__a22o_1
XU$$462 U$$462/A U$$498/B VGND VGND VPWR VPWR U$$462/X sky130_fd_sc_hd__xor2_1
XU$$473 U$$882/B1 U$$479/A2 U$$747/B1 U$$479/B2 VGND VGND VPWR VPWR U$$474/A sky130_fd_sc_hd__a22o_1
XU$$484 U$$484/A U$$504/B VGND VGND VPWR VPWR U$$484/X sky130_fd_sc_hd__xor2_1
XU$$495 U$$632/A1 U$$497/A2 U$$632/B1 U$$497/B2 VGND VGND VPWR VPWR U$$496/A sky130_fd_sc_hd__a22o_1
XFILLER_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_94_3 U$$3919/X U$$4052/X U$$4185/X VGND VGND VPWR VPWR dadda_fa_3_95_1/B
+ dadda_fa_3_94_3/B sky130_fd_sc_hd__fa_1
XFILLER_145_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_87_2 U$$4437/X input242/X dadda_fa_2_87_2/CIN VGND VGND VPWR VPWR dadda_fa_3_88_1/A
+ dadda_fa_3_87_3/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_64_1 dadda_fa_5_64_1/A dadda_fa_5_64_1/B dadda_fa_5_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_65_0/B dadda_fa_7_64_0/A sky130_fd_sc_hd__fa_1
XFILLER_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_57_0 dadda_fa_5_57_0/A dadda_fa_5_57_0/B dadda_fa_5_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_58_0/A dadda_fa_6_57_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_56_8 dadda_fa_1_56_8/A dadda_fa_1_56_8/B dadda_fa_1_56_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_57_3/A dadda_fa_3_56_0/A sky130_fd_sc_hd__fa_1
XFILLER_28_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_103_0 U$$2739/Y U$$2873/X U$$3006/X VGND VGND VPWR VPWR dadda_fa_3_104_2/B
+ dadda_fa_3_103_3/B sky130_fd_sc_hd__fa_1
XFILLER_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1190 U$$94/A1 U$$1194/A2 U$$96/A1 U$$1194/B2 VGND VGND VPWR VPWR U$$1191/A sky130_fd_sc_hd__a22o_1
XFILLER_149_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_82_1 U$$1634/X U$$1767/X U$$1900/X VGND VGND VPWR VPWR dadda_fa_2_83_1/CIN
+ dadda_fa_2_82_4/A sky130_fd_sc_hd__fa_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1707 fanout1708/X VGND VGND VPWR VPWR U$$4353/A1 sky130_fd_sc_hd__buf_4
XFILLER_172_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1718 input107/X VGND VGND VPWR VPWR fanout1718/X sky130_fd_sc_hd__buf_4
Xfanout720 U$$3912/B2 VGND VGND VPWR VPWR U$$3906/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_75_0 U$$1620/X U$$1753/X U$$1886/X VGND VGND VPWR VPWR dadda_fa_2_76_0/B
+ dadda_fa_2_75_3/B sky130_fd_sc_hd__fa_1
XFILLER_131_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1729 input105/X VGND VGND VPWR VPWR U$$922/A1 sky130_fd_sc_hd__buf_6
Xfanout731 U$$3704/X VGND VGND VPWR VPWR U$$3791/B2 sky130_fd_sc_hd__buf_6
XFILLER_120_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout742 U$$3567/X VGND VGND VPWR VPWR U$$3658/B2 sky130_fd_sc_hd__buf_4
Xfanout753 U$$3293/X VGND VGND VPWR VPWR U$$3340/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout764 U$$3156/X VGND VGND VPWR VPWR U$$3245/B2 sky130_fd_sc_hd__buf_2
Xfanout775 U$$3019/X VGND VGND VPWR VPWR U$$3122/B2 sky130_fd_sc_hd__clkbuf_2
Xfanout786 U$$2882/X VGND VGND VPWR VPWR U$$3011/B2 sky130_fd_sc_hd__buf_4
Xfanout797 U$$2844/B2 VGND VGND VPWR VPWR U$$2804/B2 sky130_fd_sc_hd__buf_4
XFILLER_100_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3509 U$$3509/A1 U$$3511/A2 U$$3509/B1 U$$3511/B2 VGND VGND VPWR VPWR U$$3510/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2808 U$$4315/A1 U$$2874/A2 U$$4454/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2809/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2819 U$$2819/A U$$2871/B VGND VGND VPWR VPWR U$$2819/X sky130_fd_sc_hd__xor2_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_422_ _422_/CLK _422_/D VGND VGND VPWR VPWR _422_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_353_ _353_/CLK _353_/D VGND VGND VPWR VPWR _353_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_284_ _416_/CLK _284_/D VGND VGND VPWR VPWR _284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_97_1 dadda_fa_3_97_1/A dadda_fa_3_97_1/B dadda_fa_3_97_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_0/CIN dadda_fa_4_97_2/A sky130_fd_sc_hd__fa_1
XFILLER_6_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_74_0 dadda_fa_6_74_0/A dadda_fa_6_74_0/B dadda_fa_6_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_75_0/B dadda_fa_7_74_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_170_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 a[16] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_119_0 U$$3835/Y U$$3969/X U$$4102/X VGND VGND VPWR VPWR dadda_fa_5_120_0/CIN
+ dadda_fa_5_119_1/B sky130_fd_sc_hd__fa_1
XFILLER_80_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$270 U$$270/A U$$274/A VGND VGND VPWR VPWR U$$270/X sky130_fd_sc_hd__xor2_1
XU$$281 U$$281/A U$$313/B VGND VGND VPWR VPWR U$$281/X sky130_fd_sc_hd__xor2_1
XU$$292 U$$18/A1 U$$312/A2 U$$20/A1 U$$312/B2 VGND VGND VPWR VPWR U$$293/A sky130_fd_sc_hd__a22o_1
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$819_1913 VGND VGND VPWR VPWR U$$819_1913/HI U$$819/B1 sky130_fd_sc_hd__conb_1
XFILLER_158_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$6 _302_/Q _174_/Q VGND VGND VPWR VPWR final_adder.U$$6/COUT final_adder.U$$6/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_161_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput301 output301/A VGND VGND VPWR VPWR o[24] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_0 U$$2984/X U$$3117/X U$$3250/X VGND VGND VPWR VPWR dadda_fa_3_93_0/B
+ dadda_fa_3_92_2/B sky130_fd_sc_hd__fa_1
Xoutput312 output312/A VGND VGND VPWR VPWR o[34] sky130_fd_sc_hd__buf_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput323 output323/A VGND VGND VPWR VPWR o[44] sky130_fd_sc_hd__buf_2
Xoutput334 output334/A VGND VGND VPWR VPWR o[54] sky130_fd_sc_hd__buf_2
Xoutput345 output345/A VGND VGND VPWR VPWR o[64] sky130_fd_sc_hd__buf_2
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput356 output356/A VGND VGND VPWR VPWR o[74] sky130_fd_sc_hd__buf_2
Xoutput367 output367/A VGND VGND VPWR VPWR o[84] sky130_fd_sc_hd__buf_2
Xoutput378 output378/A VGND VGND VPWR VPWR o[94] sky130_fd_sc_hd__buf_2
Xdadda_ha_4_118_2 U$$4499/X input149/X VGND VGND VPWR VPWR dadda_fa_5_119_1/A dadda_ha_4_118_2/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_142_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_6 dadda_fa_1_61_6/A dadda_fa_1_61_6/B dadda_fa_1_61_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_62_2/B dadda_fa_2_61_5/B sky130_fd_sc_hd__fa_1
XFILLER_56_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_5 U$$2775/X U$$2908/X U$$3041/X VGND VGND VPWR VPWR dadda_fa_2_55_2/A
+ dadda_fa_2_54_5/A sky130_fd_sc_hd__fa_1
XFILLER_83_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_47_4 U$$1697/X U$$1830/X U$$1963/X VGND VGND VPWR VPWR dadda_fa_2_48_2/CIN
+ dadda_fa_2_47_5/B sky130_fd_sc_hd__fa_1
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_17_2 dadda_fa_4_17_2/A dadda_fa_4_17_2/B dadda_ha_3_17_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_18_0/CIN dadda_fa_5_17_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_23_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_91_0 dadda_fa_7_91_0/A dadda_fa_7_91_0/B dadda_fa_7_91_0/CIN VGND VGND
+ VPWR VPWR _388_/D _259_/D sky130_fd_sc_hd__fa_1
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1504 U$$1491/B VGND VGND VPWR VPWR U$$1475/B sky130_fd_sc_hd__buf_6
Xfanout1515 U$$981/B1 VGND VGND VPWR VPWR U$$2762/B1 sky130_fd_sc_hd__clkbuf_2
Xfanout1526 input126/X VGND VGND VPWR VPWR U$$981/A1 sky130_fd_sc_hd__buf_6
Xfanout1537 U$$3580/B1 VGND VGND VPWR VPWR U$$840/B1 sky130_fd_sc_hd__buf_4
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout550 U$$2733/A2 VGND VGND VPWR VPWR U$$2737/A2 sky130_fd_sc_hd__buf_4
Xfanout1548 U$$4516/A1 VGND VGND VPWR VPWR U$$678/B1 sky130_fd_sc_hd__buf_2
Xfanout561 U$$2470/X VGND VGND VPWR VPWR fanout561/X sky130_fd_sc_hd__clkbuf_16
XU$$4007 U$$4416/B1 U$$4057/A2 U$$4283/A1 U$$4057/B2 VGND VGND VPWR VPWR U$$4008/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1559 U$$3966/A1 VGND VGND VPWR VPWR U$$4375/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout572 U$$2282/A2 VGND VGND VPWR VPWR U$$2252/A2 sky130_fd_sc_hd__buf_6
XU$$4018 U$$4018/A U$$4098/B VGND VGND VPWR VPWR U$$4018/X sky130_fd_sc_hd__xor2_1
Xfanout583 U$$2181/A2 VGND VGND VPWR VPWR U$$2189/A2 sky130_fd_sc_hd__buf_6
XU$$4029 U$$4440/A1 U$$4045/A2 U$$4440/B1 U$$4045/B2 VGND VGND VPWR VPWR U$$4030/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_924 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout594 U$$1859/A2 VGND VGND VPWR VPWR U$$1829/A2 sky130_fd_sc_hd__buf_4
XFILLER_46_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3306 U$$3580/A1 U$$3306/A2 U$$3580/B1 U$$3306/B2 VGND VGND VPWR VPWR U$$3307/A
+ sky130_fd_sc_hd__a22o_1
XU$$3317 U$$3317/A U$$3341/B VGND VGND VPWR VPWR U$$3317/X sky130_fd_sc_hd__xor2_1
XU$$3328 U$$4287/A1 U$$3338/A2 U$$4426/A1 U$$3338/B2 VGND VGND VPWR VPWR U$$3329/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3339 U$$3339/A U$$3341/B VGND VGND VPWR VPWR U$$3339/X sky130_fd_sc_hd__xor2_1
XU$$4487_1891 VGND VGND VPWR VPWR U$$4487_1891/HI U$$4487/B sky130_fd_sc_hd__conb_1
XU$$2605 U$$2740/A VGND VGND VPWR VPWR U$$2605/Y sky130_fd_sc_hd__inv_1
XU$$2616 U$$2616/A U$$2668/B VGND VGND VPWR VPWR U$$2616/X sky130_fd_sc_hd__xor2_1
XU$$2627 U$$2762/B1 U$$2665/A2 U$$2629/A1 U$$2665/B2 VGND VGND VPWR VPWR U$$2628/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2638 U$$2638/A U$$2678/B VGND VGND VPWR VPWR U$$2638/X sky130_fd_sc_hd__xor2_1
XU$$1904 U$$1904/A U$$1910/B VGND VGND VPWR VPWR U$$1904/X sky130_fd_sc_hd__xor2_1
XFILLER_62_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2649 U$$183/A1 U$$2681/A2 U$$870/A1 U$$2681/B2 VGND VGND VPWR VPWR U$$2650/A sky130_fd_sc_hd__a22o_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1915 U$$4107/A1 U$$1915/A2 U$$1915/B1 U$$1915/B2 VGND VGND VPWR VPWR U$$1916/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1926 U$$3022/A1 U$$1964/A2 U$$3022/B1 U$$1964/B2 VGND VGND VPWR VPWR U$$1927/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1937 U$$1937/A U$$1971/B VGND VGND VPWR VPWR U$$1937/X sky130_fd_sc_hd__xor2_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1948 U$$2631/B1 U$$2006/A2 U$$852/B1 U$$2006/B2 VGND VGND VPWR VPWR U$$1949/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1959 U$$1959/A U$$1963/B VGND VGND VPWR VPWR U$$1959/X sky130_fd_sc_hd__xor2_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_405_ _405_/CLK _405_/D VGND VGND VPWR VPWR _405_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_336_ _344_/CLK _336_/D VGND VGND VPWR VPWR _336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_267_ _397_/CLK _267_/D VGND VGND VPWR VPWR _267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_198_ _344_/CLK _198_/D VGND VGND VPWR VPWR _198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_71_5 dadda_fa_2_71_5/A dadda_fa_2_71_5/B dadda_fa_2_71_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_2/A dadda_fa_4_71_0/A sky130_fd_sc_hd__fa_1
XFILLER_111_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_64_4 dadda_fa_2_64_4/A dadda_fa_2_64_4/B dadda_fa_2_64_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_1/CIN dadda_fa_3_64_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_57_3 dadda_fa_2_57_3/A dadda_fa_2_57_3/B dadda_fa_2_57_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_1/B dadda_fa_3_57_3/B sky130_fd_sc_hd__fa_1
XFILLER_77_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$11 U$$11/A U$$9/B VGND VGND VPWR VPWR U$$11/X sky130_fd_sc_hd__xor2_1
XU$$22 U$$22/A1 U$$8/A2 U$$24/A1 U$$8/B2 VGND VGND VPWR VPWR U$$23/A sky130_fd_sc_hd__a22o_1
XU$$33 U$$33/A U$$49/B VGND VGND VPWR VPWR U$$33/X sky130_fd_sc_hd__xor2_1
XU$$44 U$$44/A1 U$$48/A2 U$$46/A1 U$$48/B2 VGND VGND VPWR VPWR U$$45/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_27_1 dadda_fa_5_27_1/A dadda_fa_5_27_1/B dadda_fa_5_27_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_28_0/B dadda_fa_7_27_0/A sky130_fd_sc_hd__fa_2
XU$$55 U$$55/A U$$87/B VGND VGND VPWR VPWR U$$55/X sky130_fd_sc_hd__xor2_1
XU$$3840 U$$3838/Y input52/X U$$3836/A U$$3839/X U$$3836/Y VGND VGND VPWR VPWR U$$3840/X
+ sky130_fd_sc_hd__a32o_2
XU$$66 U$$66/A1 U$$96/A2 U$$66/B1 U$$96/B2 VGND VGND VPWR VPWR U$$67/A sky130_fd_sc_hd__a22o_1
XU$$3851 U$$3851/A U$$3867/B VGND VGND VPWR VPWR U$$3851/X sky130_fd_sc_hd__xor2_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3862 U$$3999/A1 U$$3872/A2 U$$3999/B1 U$$3872/B2 VGND VGND VPWR VPWR U$$3863/A
+ sky130_fd_sc_hd__a22o_1
XU$$3873 U$$3873/A U$$3893/B VGND VGND VPWR VPWR U$$3873/X sky130_fd_sc_hd__xor2_1
XU$$77 U$$77/A U$$77/B VGND VGND VPWR VPWR U$$77/X sky130_fd_sc_hd__xor2_1
XFILLER_18_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$88 U$$88/A1 U$$96/A2 U$$88/B1 U$$96/B2 VGND VGND VPWR VPWR U$$89/A sky130_fd_sc_hd__a22o_1
XU$$99 U$$99/A U$$99/B VGND VGND VPWR VPWR U$$99/X sky130_fd_sc_hd__xor2_1
XU$$3884 U$$3884/A1 U$$3970/A2 U$$4434/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3885/A
+ sky130_fd_sc_hd__a22o_1
XU$$3895 U$$3895/A U$$3907/B VGND VGND VPWR VPWR U$$3895/X sky130_fd_sc_hd__xor2_1
XFILLER_36_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_101_1 dadda_fa_5_101_1/A dadda_fa_5_101_1/B dadda_fa_5_101_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_102_0/B dadda_fa_7_101_0/A sky130_fd_sc_hd__fa_1
XFILLER_173_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_835 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_39_2 U$$883/X U$$1016/X VGND VGND VPWR VPWR dadda_fa_2_40_4/CIN dadda_fa_3_39_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_102_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_924 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_52_2 U$$1175/X U$$1308/X U$$1441/X VGND VGND VPWR VPWR dadda_fa_2_53_1/A
+ dadda_fa_2_52_4/A sky130_fd_sc_hd__fa_1
XFILLER_28_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_45_1 U$$496/X U$$629/X U$$762/X VGND VGND VPWR VPWR dadda_fa_2_46_2/B
+ dadda_fa_2_45_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_22_0 dadda_fa_4_22_0/A dadda_fa_4_22_0/B dadda_fa_4_22_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_23_0/A dadda_fa_5_22_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_38_0 U$$83/X U$$216/X U$$349/X VGND VGND VPWR VPWR dadda_fa_2_39_4/B dadda_fa_2_38_5/B
+ sky130_fd_sc_hd__fa_1
XFILLER_169_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1005 final_adder.U$$234/A final_adder.U$$735/X final_adder.U$$235/A2
+ VGND VGND VPWR VPWR final_adder.U$$1045/B sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$1027 final_adder.U$$3/SUM final_adder.U$$1027/B VGND VGND VPWR VPWR
+ output318/A sky130_fd_sc_hd__xor2_1
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1038 final_adder.U$$240/A final_adder.U$$621/X VGND VGND VPWR VPWR
+ output290/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1049 final_adder.U$$230/B final_adder.U$$1049/B VGND VGND VPWR VPWR
+ output302/A sky130_fd_sc_hd__xor2_1
XFILLER_164_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_74_3 dadda_fa_3_74_3/A dadda_fa_3_74_3/B dadda_fa_3_74_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_1/B dadda_fa_4_74_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1301 fanout1309/X VGND VGND VPWR VPWR U$$3893/B sky130_fd_sc_hd__buf_4
Xdadda_fa_3_67_2 dadda_fa_3_67_2/A dadda_fa_3_67_2/B dadda_fa_3_67_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_1/A dadda_fa_4_67_2/B sky130_fd_sc_hd__fa_1
Xfanout1312 U$$3740/B VGND VGND VPWR VPWR U$$3836/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1323 U$$913/B VGND VGND VPWR VPWR U$$875/B sky130_fd_sc_hd__buf_6
Xfanout1334 U$$3698/A VGND VGND VPWR VPWR U$$3681/B sky130_fd_sc_hd__buf_6
Xfanout1345 input47/X VGND VGND VPWR VPWR U$$3524/B sky130_fd_sc_hd__clkbuf_4
Xfanout1356 fanout1364/X VGND VGND VPWR VPWR U$$3208/B sky130_fd_sc_hd__buf_6
Xfanout1367 input40/X VGND VGND VPWR VPWR U$$3107/B sky130_fd_sc_hd__buf_6
Xfanout1378 U$$2990/B VGND VGND VPWR VPWR U$$2944/B sky130_fd_sc_hd__buf_6
Xfanout391 U$$963/X VGND VGND VPWR VPWR U$$1087/A2 sky130_fd_sc_hd__buf_6
Xfanout1389 U$$2873/B VGND VGND VPWR VPWR U$$2876/A sky130_fd_sc_hd__buf_8
Xdadda_fa_6_37_0 dadda_fa_6_37_0/A dadda_fa_6_37_0/B dadda_fa_6_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_38_0/B dadda_fa_7_37_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_19_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3103 U$$3103/A U$$3107/B VGND VGND VPWR VPWR U$$3103/X sky130_fd_sc_hd__xor2_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3114 U$$3249/B1 U$$3118/A2 U$$4486/A1 U$$3118/B2 VGND VGND VPWR VPWR U$$3115/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3125 U$$3125/A U$$3150/A VGND VGND VPWR VPWR U$$3125/X sky130_fd_sc_hd__xor2_1
XU$$3136 U$$4093/B1 U$$3148/A2 U$$3684/B1 U$$3148/B2 VGND VGND VPWR VPWR U$$3137/A
+ sky130_fd_sc_hd__a22o_1
XU$$2402 U$$2402/A U$$2402/B VGND VGND VPWR VPWR U$$2402/X sky130_fd_sc_hd__xor2_1
XU$$3147 U$$3147/A U$$3147/B VGND VGND VPWR VPWR U$$3147/X sky130_fd_sc_hd__xor2_1
XU$$2413 U$$3920/A1 U$$2413/A2 U$$908/A1 U$$2413/B2 VGND VGND VPWR VPWR U$$2414/A
+ sky130_fd_sc_hd__a22o_1
XU$$3158 U$$3158/A U$$3196/B VGND VGND VPWR VPWR U$$3158/X sky130_fd_sc_hd__xor2_1
XFILLER_74_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2424 U$$2424/A U$$2456/B VGND VGND VPWR VPWR U$$2424/X sky130_fd_sc_hd__xor2_1
XU$$3169 U$$566/A1 U$$3257/A2 U$$979/A1 U$$3257/B2 VGND VGND VPWR VPWR U$$3170/A sky130_fd_sc_hd__a22o_1
XU$$2435 U$$2707/B1 U$$2443/A2 U$$2574/A1 U$$2443/B2 VGND VGND VPWR VPWR U$$2436/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1701 U$$1701/A U$$1703/B VGND VGND VPWR VPWR U$$1701/X sky130_fd_sc_hd__xor2_1
XU$$2446 U$$2446/A U$$2446/B VGND VGND VPWR VPWR U$$2446/X sky130_fd_sc_hd__xor2_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1712 U$$479/A1 U$$1720/A2 U$$479/B1 U$$1720/B2 VGND VGND VPWR VPWR U$$1713/A sky130_fd_sc_hd__a22o_1
XU$$2457 U$$950/A1 U$$2459/A2 U$$952/A1 U$$2459/B2 VGND VGND VPWR VPWR U$$2458/A sky130_fd_sc_hd__a22o_1
XU$$2468 U$$2575/B VGND VGND VPWR VPWR U$$2468/Y sky130_fd_sc_hd__inv_1
XU$$1723 U$$1723/A U$$1727/B VGND VGND VPWR VPWR U$$1723/X sky130_fd_sc_hd__xor2_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1734 U$$3376/B1 U$$1774/A2 U$$3243/A1 U$$1774/B2 VGND VGND VPWR VPWR U$$1735/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2479 U$$2479/A U$$2545/B VGND VGND VPWR VPWR U$$2479/X sky130_fd_sc_hd__xor2_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1745 U$$1745/A U$$1761/B VGND VGND VPWR VPWR U$$1745/X sky130_fd_sc_hd__xor2_1
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1756 U$$521/B1 U$$1758/A2 U$$386/B1 U$$1758/B2 VGND VGND VPWR VPWR U$$1757/A sky130_fd_sc_hd__a22o_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1767 U$$1767/A U$$1777/B VGND VGND VPWR VPWR U$$1767/X sky130_fd_sc_hd__xor2_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1778 U$$4244/A1 U$$1778/A2 U$$1778/B1 U$$1778/B2 VGND VGND VPWR VPWR U$$1779/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1789 U$$3022/A1 U$$1829/A2 U$$3022/B1 U$$1829/B2 VGND VGND VPWR VPWR U$$1790/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_319_ _319_/CLK _319_/D VGND VGND VPWR VPWR _319_/Q sky130_fd_sc_hd__dfxtp_1
Xinput11 a[19] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput22 a[29] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_1
Xinput33 a[39] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
Xinput44 a[49] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__buf_4
Xinput55 a[59] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__clkbuf_1
Xinput66 b[10] VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__clkbuf_4
Xinput77 b[20] VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput88 b[30] VGND VGND VPWR VPWR input88/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput99 b[40] VGND VGND VPWR VPWR input99/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4_1829 VGND VGND VPWR VPWR U$$4_1829/HI U$$4/A3 sky130_fd_sc_hd__conb_1
Xdadda_fa_2_62_1 dadda_fa_2_62_1/A dadda_fa_2_62_1/B dadda_fa_2_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_0/CIN dadda_fa_3_62_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$408 final_adder.U$$412/B final_adder.U$$408/B VGND VGND VPWR VPWR
+ final_adder.U$$532/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$419 final_adder.U$$418/B final_adder.U$$297/X final_adder.U$$293/X
+ VGND VGND VPWR VPWR final_adder.U$$419/X sky130_fd_sc_hd__a21o_1
XFILLER_85_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_55_0 dadda_fa_2_55_0/A dadda_fa_2_55_0/B dadda_fa_2_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_0/B dadda_fa_3_55_2/B sky130_fd_sc_hd__fa_1
XFILLER_84_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4360 U$$4360/A U$$4360/B VGND VGND VPWR VPWR U$$4360/X sky130_fd_sc_hd__xor2_1
XU$$4371 U$$4508/A1 U$$4373/A2 U$$4508/B1 U$$4373/B2 VGND VGND VPWR VPWR U$$4372/A
+ sky130_fd_sc_hd__a22o_1
XU$$4382 U$$4382/A U$$4383/A VGND VGND VPWR VPWR U$$4382/X sky130_fd_sc_hd__xor2_1
XU$$4393 U$$4393/A U$$4393/B VGND VGND VPWR VPWR U$$4393/X sky130_fd_sc_hd__xor2_1
XU$$3670 U$$4492/A1 U$$3692/A2 U$$4492/B1 U$$3692/B2 VGND VGND VPWR VPWR U$$3671/A
+ sky130_fd_sc_hd__a22o_1
XU$$3681 U$$3681/A U$$3681/B VGND VGND VPWR VPWR U$$3681/X sky130_fd_sc_hd__xor2_1
XU$$3692 U$$3692/A1 U$$3692/A2 U$$3692/B1 U$$3692/B2 VGND VGND VPWR VPWR U$$3693/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_9_0 U$$291/X U$$424/X U$$557/X VGND VGND VPWR VPWR dadda_fa_6_10_0/A dadda_fa_6_9_0/CIN
+ sky130_fd_sc_hd__fa_1
XU$$2980 U$$2980/A U$$3014/A VGND VGND VPWR VPWR U$$2980/X sky130_fd_sc_hd__xor2_1
XFILLER_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2991 U$$251/A1 U$$2991/A2 U$$251/B1 U$$2991/B2 VGND VGND VPWR VPWR U$$2992/A sky130_fd_sc_hd__a22o_1
XFILLER_34_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_84_2 dadda_fa_4_84_2/A dadda_fa_4_84_2/B dadda_fa_4_84_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_85_0/CIN dadda_fa_5_84_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_77_1 dadda_fa_4_77_1/A dadda_fa_4_77_1/B dadda_fa_4_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_78_0/B dadda_fa_5_77_1/B sky130_fd_sc_hd__fa_1
XFILLER_134_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_54_0 dadda_fa_7_54_0/A dadda_fa_7_54_0/B dadda_fa_7_54_0/CIN VGND VGND
+ VPWR VPWR _351_/D _222_/D sky130_fd_sc_hd__fa_1
XFILLER_103_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$931 final_adder.U$$160/A final_adder.U$$869/X final_adder.U$$931/B1
+ VGND VGND VPWR VPWR final_adder.U$$931/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$953 final_adder.U$$182/A final_adder.U$$891/X final_adder.U$$953/B1
+ VGND VGND VPWR VPWR final_adder.U$$953/X sky130_fd_sc_hd__a21o_1
XFILLER_29_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$803 U$$803/A1 U$$809/A2 U$$805/A1 U$$809/B2 VGND VGND VPWR VPWR U$$804/A sky130_fd_sc_hd__a22o_1
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$975 final_adder.U$$204/A final_adder.U$$817/X final_adder.U$$975/B1
+ VGND VGND VPWR VPWR final_adder.U$$975/X sky130_fd_sc_hd__a21o_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$814 U$$814/A U$$820/B VGND VGND VPWR VPWR U$$814/X sky130_fd_sc_hd__xor2_1
XU$$825 U$$959/A U$$825/B VGND VGND VPWR VPWR U$$825/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$997 final_adder.U$$226/A final_adder.U$$727/X final_adder.U$$997/B1
+ VGND VGND VPWR VPWR final_adder.U$$997/X sky130_fd_sc_hd__a21o_1
XFILLER_84_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$836 U$$973/A1 U$$904/A2 U$$973/B1 U$$904/B2 VGND VGND VPWR VPWR U$$837/A sky130_fd_sc_hd__a22o_1
XFILLER_73_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$847 U$$847/A U$$875/B VGND VGND VPWR VPWR U$$847/X sky130_fd_sc_hd__xor2_1
XU$$858 U$$995/A1 U$$898/A2 U$$997/A1 U$$898/B2 VGND VGND VPWR VPWR U$$859/A sky130_fd_sc_hd__a22o_1
XFILLER_44_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1008 U$$1008/A U$$980/B VGND VGND VPWR VPWR U$$1008/X sky130_fd_sc_hd__xor2_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$869 U$$869/A U$$925/B VGND VGND VPWR VPWR U$$869/X sky130_fd_sc_hd__xor2_1
XU$$1019 U$$60/A1 U$$999/A2 U$$62/A1 U$$999/B2 VGND VGND VPWR VPWR U$$1020/A sky130_fd_sc_hd__a22o_1
XFILLER_71_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_72_0 dadda_fa_3_72_0/A dadda_fa_3_72_0/B dadda_fa_3_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_0/B dadda_fa_4_72_1/CIN sky130_fd_sc_hd__fa_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1120 U$$3610/B1 VGND VGND VPWR VPWR U$$3338/A1 sky130_fd_sc_hd__buf_4
Xfanout1131 U$$4432/A1 VGND VGND VPWR VPWR U$$4158/A1 sky130_fd_sc_hd__buf_6
Xfanout1142 U$$2923/A1 VGND VGND VPWR VPWR U$$729/B1 sky130_fd_sc_hd__buf_4
XFILLER_26_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1153 U$$4291/A1 VGND VGND VPWR VPWR U$$4428/A1 sky130_fd_sc_hd__buf_6
Xfanout1164 U$$40/B1 VGND VGND VPWR VPWR U$$2780/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1175 U$$4424/A1 VGND VGND VPWR VPWR U$$4150/A1 sky130_fd_sc_hd__buf_6
Xfanout1186 U$$3870/B1 VGND VGND VPWR VPWR U$$3322/B1 sky130_fd_sc_hd__buf_6
XFILLER_94_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1197 U$$982/B VGND VGND VPWR VPWR U$$980/B sky130_fd_sc_hd__buf_6
XFILLER_47_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2210 U$$840/A1 U$$2252/A2 U$$840/B1 U$$2252/B2 VGND VGND VPWR VPWR U$$2211/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_101_0 dadda_fa_4_101_0/A dadda_fa_4_101_0/B dadda_fa_4_101_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_102_0/A dadda_fa_5_101_1/A sky130_fd_sc_hd__fa_1
XU$$2221 U$$2221/A U$$2231/B VGND VGND VPWR VPWR U$$2221/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_34_5 U$$2336/X U$$2412/B input184/X VGND VGND VPWR VPWR dadda_fa_3_35_2/A
+ dadda_fa_4_34_0/A sky130_fd_sc_hd__fa_2
XU$$2232 U$$999/A1 U$$2272/A2 U$$999/B1 U$$2272/B2 VGND VGND VPWR VPWR U$$2233/A sky130_fd_sc_hd__a22o_1
XU$$2243 U$$2243/A U$$2249/B VGND VGND VPWR VPWR U$$2243/X sky130_fd_sc_hd__xor2_1
XU$$2254 U$$2665/A1 U$$2254/A2 U$$2665/B1 U$$2254/B2 VGND VGND VPWR VPWR U$$2255/A
+ sky130_fd_sc_hd__a22o_1
XU$$2265 U$$2265/A U$$2269/B VGND VGND VPWR VPWR U$$2265/X sky130_fd_sc_hd__xor2_1
XU$$1520 U$$1520/A U$$1568/B VGND VGND VPWR VPWR U$$1520/X sky130_fd_sc_hd__xor2_1
XFILLER_16_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1531 U$$983/A1 U$$1567/A2 U$$983/B1 U$$1567/B2 VGND VGND VPWR VPWR U$$1532/A sky130_fd_sc_hd__a22o_1
XU$$2276 U$$4468/A1 U$$2326/A2 U$$4470/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2277/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1542 U$$1542/A U$$1570/B VGND VGND VPWR VPWR U$$1542/X sky130_fd_sc_hd__xor2_1
XU$$2287 U$$2287/A U$$2327/B VGND VGND VPWR VPWR U$$2287/X sky130_fd_sc_hd__xor2_1
XU$$1553 U$$729/B1 U$$1563/A2 U$$596/A1 U$$1563/B2 VGND VGND VPWR VPWR U$$1554/A sky130_fd_sc_hd__a22o_1
XFILLER_16_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2298 U$$2707/B1 U$$2310/A2 U$$2574/A1 U$$2310/B2 VGND VGND VPWR VPWR U$$2299/A
+ sky130_fd_sc_hd__a22o_1
XU$$1564 U$$1564/A U$$1564/B VGND VGND VPWR VPWR U$$1564/X sky130_fd_sc_hd__xor2_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1575 U$$616/A1 U$$1575/A2 U$$481/A1 U$$1575/B2 VGND VGND VPWR VPWR U$$1576/A sky130_fd_sc_hd__a22o_1
XU$$1586 U$$1586/A U$$1618/B VGND VGND VPWR VPWR U$$1586/X sky130_fd_sc_hd__xor2_1
XFILLER_33_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1597 U$$3239/B1 U$$1641/A2 U$$3106/A1 U$$1641/B2 VGND VGND VPWR VPWR U$$1598/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_94_1 dadda_fa_5_94_1/A dadda_fa_5_94_1/B dadda_fa_5_94_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_95_0/B dadda_fa_7_94_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_87_0 dadda_fa_5_87_0/A dadda_fa_5_87_0/B dadda_fa_5_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_88_0/A dadda_fa_6_87_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_79_7 U$$3889/X U$$4022/X U$$4155/X VGND VGND VPWR VPWR dadda_fa_2_80_2/CIN
+ dadda_fa_2_79_5/CIN sky130_fd_sc_hd__fa_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$205 final_adder.U$$204/B final_adder.U$$975/B1 final_adder.U$$205/B1
+ VGND VGND VPWR VPWR final_adder.U$$205/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$216 final_adder.U$$216/A final_adder.U$$216/B VGND VGND VPWR VPWR
+ final_adder.U$$344/B sky130_fd_sc_hd__and2_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$227 final_adder.U$$226/B final_adder.U$$997/B1 final_adder.U$$227/B1
+ VGND VGND VPWR VPWR final_adder.U$$227/X sky130_fd_sc_hd__a21o_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$238 final_adder.U$$238/A final_adder.U$$238/B VGND VGND VPWR VPWR
+ final_adder.U$$366/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$249 final_adder.U$$7/SUM final_adder.U$$6/COUT final_adder.U$$7/COUT
+ VGND VGND VPWR VPWR final_adder.U$$249/X sky130_fd_sc_hd__a21o_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4190 U$$4464/A1 U$$4190/A2 U$$4464/B1 U$$4190/B2 VGND VGND VPWR VPWR U$$4191/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_103_2 dadda_fa_3_103_2/A dadda_fa_3_103_2/B dadda_fa_3_103_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_104_1/A dadda_fa_4_103_2/B sky130_fd_sc_hd__fa_1
XFILLER_150_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput201 c[4] VGND VGND VPWR VPWR input201/X sky130_fd_sc_hd__clkbuf_4
XFILLER_89_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput212 c[5] VGND VGND VPWR VPWR input212/X sky130_fd_sc_hd__clkbuf_4
XFILLER_88_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput223 c[6] VGND VGND VPWR VPWR input223/X sky130_fd_sc_hd__clkbuf_4
Xinput234 c[7] VGND VGND VPWR VPWR input234/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput245 c[8] VGND VGND VPWR VPWR input245/X sky130_fd_sc_hd__clkbuf_4
XFILLER_102_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput256 c[9] VGND VGND VPWR VPWR input256/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_0_67_5 U$$2136/X U$$2269/X U$$2402/X VGND VGND VPWR VPWR dadda_fa_1_68_7/A
+ dadda_fa_2_67_0/A sky130_fd_sc_hd__fa_1
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_117_0 dadda_fa_6_117_0/A dadda_fa_6_117_0/B dadda_fa_6_117_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_118_0/B dadda_fa_7_117_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_124_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$750 final_adder.U$$782/B final_adder.U$$750/B VGND VGND VPWR VPWR
+ final_adder.U$$750/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$761 final_adder.U$$760/B final_adder.U$$681/X final_adder.U$$649/X
+ VGND VGND VPWR VPWR final_adder.U$$761/X sky130_fd_sc_hd__a21o_1
XU$$600 U$$52/A1 U$$636/A2 U$$54/A1 U$$636/B2 VGND VGND VPWR VPWR U$$601/A sky130_fd_sc_hd__a22o_1
XFILLER_63_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$772 final_adder.U$$772/A final_adder.U$$772/B VGND VGND VPWR VPWR
+ final_adder.U$$772/X sky130_fd_sc_hd__and2_1
XU$$611 U$$611/A U$$643/B VGND VGND VPWR VPWR U$$611/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$783 final_adder.U$$782/B final_adder.U$$703/X final_adder.U$$671/X
+ VGND VGND VPWR VPWR final_adder.U$$783/X sky130_fd_sc_hd__a21o_1
XU$$622 U$$896/A1 U$$630/A2 U$$898/A1 U$$630/B2 VGND VGND VPWR VPWR U$$623/A sky130_fd_sc_hd__a22o_1
XFILLER_75_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_37_3 dadda_fa_3_37_3/A dadda_fa_3_37_3/B dadda_fa_3_37_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_1/B dadda_fa_4_37_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_90_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$794 final_adder.U$$794/A final_adder.U$$794/B VGND VGND VPWR VPWR
+ final_adder.U$$794/X sky130_fd_sc_hd__and2_1
XU$$633 U$$633/A U$$669/B VGND VGND VPWR VPWR U$$633/X sky130_fd_sc_hd__xor2_1
XU$$644 U$$781/A1 U$$682/A2 U$$783/A1 U$$682/B2 VGND VGND VPWR VPWR U$$645/A sky130_fd_sc_hd__a22o_1
XFILLER_17_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$655 U$$655/A U$$684/A VGND VGND VPWR VPWR U$$655/X sky130_fd_sc_hd__xor2_1
XU$$666 U$$803/A1 U$$674/A2 U$$805/A1 U$$674/B2 VGND VGND VPWR VPWR U$$667/A sky130_fd_sc_hd__a22o_1
XU$$677 U$$677/A U$$685/A VGND VGND VPWR VPWR U$$677/X sky130_fd_sc_hd__xor2_1
XU$$688 U$$804/B U$$688/B VGND VGND VPWR VPWR U$$688/X sky130_fd_sc_hd__and2_1
XFILLER_71_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$699 U$$14/A1 U$$743/A2 U$$16/A1 U$$743/B2 VGND VGND VPWR VPWR U$$700/A sky130_fd_sc_hd__a22o_1
XFILLER_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$956_1915 VGND VGND VPWR VPWR U$$956_1915/HI U$$956/B1 sky130_fd_sc_hd__conb_1
XFILLER_13_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_32_2 U$$869/X U$$1002/X U$$1135/X VGND VGND VPWR VPWR dadda_fa_3_33_1/A
+ dadda_fa_3_32_3/A sky130_fd_sc_hd__fa_1
XFILLER_81_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2040 U$$2175/B1 U$$2044/A2 U$$2042/A1 U$$2044/B2 VGND VGND VPWR VPWR U$$2041/A
+ sky130_fd_sc_hd__a22o_1
XU$$2051 U$$2051/A U$$2053/B VGND VGND VPWR VPWR U$$2051/X sky130_fd_sc_hd__xor2_1
XU$$2062 U$$2062/A U$$2096/B VGND VGND VPWR VPWR U$$2062/X sky130_fd_sc_hd__xor2_1
XU$$2073 U$$566/A1 U$$2147/A2 U$$979/A1 U$$2147/B2 VGND VGND VPWR VPWR U$$2074/A sky130_fd_sc_hd__a22o_1
XU$$2084 U$$2084/A U$$2130/B VGND VGND VPWR VPWR U$$2084/X sky130_fd_sc_hd__xor2_1
XU$$2095 U$$3189/B1 U$$2097/A2 U$$3056/A1 U$$2097/B2 VGND VGND VPWR VPWR U$$2096/A
+ sky130_fd_sc_hd__a22o_1
XU$$1350 U$$1350/A U$$1358/B VGND VGND VPWR VPWR U$$1350/X sky130_fd_sc_hd__xor2_1
XU$$1361 U$$811/B1 U$$1361/A2 U$$678/A1 U$$1361/B2 VGND VGND VPWR VPWR U$$1362/A sky130_fd_sc_hd__a22o_1
XU$$1372 U$$1507/A VGND VGND VPWR VPWR U$$1372/Y sky130_fd_sc_hd__inv_1
XU$$1383 U$$1383/A U$$1415/B VGND VGND VPWR VPWR U$$1383/X sky130_fd_sc_hd__xor2_1
XU$$1394 U$$983/A1 U$$1426/A2 U$$983/B1 U$$1426/B2 VGND VGND VPWR VPWR U$$1395/A sky130_fd_sc_hd__a22o_1
XFILLER_148_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_84_5 U$$3367/X U$$3500/X U$$3633/X VGND VGND VPWR VPWR dadda_fa_2_85_3/CIN
+ dadda_fa_2_84_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_104_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout902 U$$1353/B2 VGND VGND VPWR VPWR U$$1359/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout913 U$$102/B2 VGND VGND VPWR VPWR U$$86/B2 sky130_fd_sc_hd__buf_4
Xfanout924 U$$4389/X VGND VGND VPWR VPWR U$$4458/B2 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_1_77_4 U$$2954/X U$$3087/X U$$3220/X VGND VGND VPWR VPWR dadda_fa_2_78_1/CIN
+ dadda_fa_2_77_4/CIN sky130_fd_sc_hd__fa_1
Xfanout935 U$$3650/A1 VGND VGND VPWR VPWR U$$4472/A1 sky130_fd_sc_hd__clkbuf_2
Xfanout946 U$$3713/A1 VGND VGND VPWR VPWR U$$973/A1 sky130_fd_sc_hd__buf_6
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout957 input97/X VGND VGND VPWR VPWR fanout957/X sky130_fd_sc_hd__buf_6
Xfanout968 fanout975/X VGND VGND VPWR VPWR U$$902/B1 sky130_fd_sc_hd__clkbuf_4
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout979 fanout984/X VGND VGND VPWR VPWR U$$3642/A1 sky130_fd_sc_hd__buf_4
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_47_2 dadda_fa_4_47_2/A dadda_fa_4_47_2/B dadda_fa_4_47_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_48_0/CIN dadda_fa_5_47_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_17_0 dadda_fa_7_17_0/A dadda_fa_7_17_0/B dadda_fa_7_17_0/CIN VGND VGND
+ VPWR VPWR _314_/D _185_/D sky130_fd_sc_hd__fa_2
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$90 _386_/Q _258_/Q VGND VGND VPWR VPWR final_adder.U$$935/B1 final_adder.U$$164/A
+ sky130_fd_sc_hd__ha_4
XFILLER_110_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_0_59_3 U$$1322/X U$$1455/X VGND VGND VPWR VPWR dadda_fa_1_60_7/B dadda_fa_2_59_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_49_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_65_2 U$$935/X U$$1068/X U$$1201/X VGND VGND VPWR VPWR dadda_fa_1_66_6/A
+ dadda_fa_1_65_8/A sky130_fd_sc_hd__fa_1
XFILLER_49_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_42_1 dadda_fa_3_42_1/A dadda_fa_3_42_1/B dadda_fa_3_42_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_0/CIN dadda_fa_4_42_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_0_58_1 U$$522/X U$$655/X U$$788/X VGND VGND VPWR VPWR dadda_fa_1_59_7/A
+ dadda_fa_1_58_8/B sky130_fd_sc_hd__fa_1
XFILLER_17_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$580 final_adder.U$$588/B final_adder.U$$580/B VGND VGND VPWR VPWR
+ final_adder.U$$700/B sky130_fd_sc_hd__and2_1
Xdadda_fa_3_35_0 dadda_fa_3_35_0/A dadda_fa_3_35_0/B dadda_fa_3_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_0/B dadda_fa_4_35_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$591 final_adder.U$$590/B final_adder.U$$475/X final_adder.U$$467/X
+ VGND VGND VPWR VPWR final_adder.U$$591/X sky130_fd_sc_hd__a21o_1
XFILLER_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$430 U$$430/A U$$480/B VGND VGND VPWR VPWR U$$430/X sky130_fd_sc_hd__xor2_1
XU$$441 U$$576/B1 U$$505/A2 U$$443/A1 U$$505/B2 VGND VGND VPWR VPWR U$$442/A sky130_fd_sc_hd__a22o_1
XU$$452 U$$452/A U$$504/B VGND VGND VPWR VPWR U$$452/X sky130_fd_sc_hd__xor2_1
XU$$463 U$$598/B1 U$$497/A2 U$$465/A1 U$$497/B2 VGND VGND VPWR VPWR U$$464/A sky130_fd_sc_hd__a22o_1
XU$$474 U$$474/A U$$480/B VGND VGND VPWR VPWR U$$474/X sky130_fd_sc_hd__xor2_1
XU$$485 U$$896/A1 U$$501/A2 U$$487/A1 U$$501/B2 VGND VGND VPWR VPWR U$$486/A sky130_fd_sc_hd__a22o_1
XU$$496 U$$496/A U$$498/B VGND VGND VPWR VPWR U$$496/X sky130_fd_sc_hd__xor2_1
XFILLER_71_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_94_4 U$$4318/X U$$4451/X input250/X VGND VGND VPWR VPWR dadda_fa_3_95_1/CIN
+ dadda_fa_3_94_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_126_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_87_3 dadda_fa_2_87_3/A dadda_fa_2_87_3/B dadda_fa_2_87_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_88_1/B dadda_fa_3_87_3/B sky130_fd_sc_hd__fa_1
XFILLER_126_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_57_1 dadda_fa_5_57_1/A dadda_fa_5_57_1/B dadda_fa_5_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_58_0/B dadda_fa_7_57_0/A sky130_fd_sc_hd__fa_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_103_1 U$$3139/X U$$3272/X U$$3405/X VGND VGND VPWR VPWR dadda_fa_3_104_2/CIN
+ dadda_fa_3_103_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1180 U$$82/B1 U$$1226/A2 U$$906/B1 U$$1226/B2 VGND VGND VPWR VPWR U$$1181/A sky130_fd_sc_hd__a22o_1
XU$$1191 U$$1191/A U$$1195/B VGND VGND VPWR VPWR U$$1191/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_124_0 dadda_fa_5_124_0/A U$$4245/X U$$4378/X VGND VGND VPWR VPWR dadda_fa_6_125_0/B
+ dadda_fa_6_124_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_148_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1006 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_82_2 U$$2033/X U$$2166/X U$$2299/X VGND VGND VPWR VPWR dadda_fa_2_83_2/A
+ dadda_fa_2_82_4/B sky130_fd_sc_hd__fa_1
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout710 U$$4043/B2 VGND VGND VPWR VPWR U$$4005/B2 sky130_fd_sc_hd__buf_2
Xfanout1708 U$$2844/B1 VGND VGND VPWR VPWR fanout1708/X sky130_fd_sc_hd__buf_4
Xfanout1719 U$$922/B1 VGND VGND VPWR VPWR U$$924/A1 sky130_fd_sc_hd__buf_6
Xfanout721 U$$3841/X VGND VGND VPWR VPWR U$$3912/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout732 U$$3833/B2 VGND VGND VPWR VPWR U$$3829/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_75_1 U$$2019/X U$$2152/X U$$2285/X VGND VGND VPWR VPWR dadda_fa_2_76_0/CIN
+ dadda_fa_2_75_3/CIN sky130_fd_sc_hd__fa_1
Xfanout743 U$$3473/B2 VGND VGND VPWR VPWR U$$3471/B2 sky130_fd_sc_hd__buf_6
XFILLER_120_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout754 U$$3378/B2 VGND VGND VPWR VPWR U$$3372/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_52_0 dadda_fa_4_52_0/A dadda_fa_4_52_0/B dadda_fa_4_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_53_0/A dadda_fa_5_52_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_68_0 U$$2537/X U$$2670/X U$$2803/X VGND VGND VPWR VPWR dadda_fa_2_69_0/B
+ dadda_fa_2_68_3/B sky130_fd_sc_hd__fa_1
XFILLER_86_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout765 U$$3257/B2 VGND VGND VPWR VPWR U$$3255/B2 sky130_fd_sc_hd__clkbuf_8
Xdadda_ha_2_102_3 U$$3802/X U$$3935/X VGND VGND VPWR VPWR dadda_fa_3_103_3/A dadda_fa_4_102_0/A
+ sky130_fd_sc_hd__ha_1
Xfanout776 U$$3118/B2 VGND VGND VPWR VPWR U$$3148/B2 sky130_fd_sc_hd__buf_4
Xfanout787 U$$279/X VGND VGND VPWR VPWR U$$362/B2 sky130_fd_sc_hd__buf_4
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout798 U$$2844/B2 VGND VGND VPWR VPWR U$$2840/B2 sky130_fd_sc_hd__buf_4
XFILLER_105_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2809 U$$2809/A U$$2876/A VGND VGND VPWR VPWR U$$2809/X sky130_fd_sc_hd__xor2_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_421_ _421_/CLK _421_/D VGND VGND VPWR VPWR _421_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ _353_/CLK _352_/D VGND VGND VPWR VPWR _352_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ _416_/CLK _283_/D VGND VGND VPWR VPWR _283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_97_2 dadda_fa_3_97_2/A dadda_fa_3_97_2/B dadda_fa_3_97_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_1/A dadda_fa_4_97_2/B sky130_fd_sc_hd__fa_1
XFILLER_127_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_67_0 dadda_fa_6_67_0/A dadda_fa_6_67_0/B dadda_fa_6_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_68_0/B dadda_fa_7_67_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_70_0 dadda_fa_0_70_0/A U$$546/X U$$679/X VGND VGND VPWR VPWR dadda_fa_1_71_6/B
+ dadda_fa_1_70_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput9 a[17] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_2
XFILLER_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_119_1 U$$4235/X U$$4368/X U$$4501/X VGND VGND VPWR VPWR dadda_fa_5_120_1/A
+ dadda_fa_5_119_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_91_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_5_6_1 U$$418/X U$$448/B VGND VGND VPWR VPWR dadda_fa_6_7_0/B dadda_fa_7_6_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_45_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$260 U$$260/A U$$260/B VGND VGND VPWR VPWR U$$260/X sky130_fd_sc_hd__xor2_1
XU$$271 U$$406/B1 U$$271/A2 U$$271/B1 U$$271/B2 VGND VGND VPWR VPWR U$$272/A sky130_fd_sc_hd__a22o_1
XFILLER_45_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$282 U$$965/B1 U$$312/A2 U$$10/A1 U$$312/B2 VGND VGND VPWR VPWR U$$283/A sky130_fd_sc_hd__a22o_1
XFILLER_32_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$293 U$$293/A U$$313/B VGND VGND VPWR VPWR U$$293/X sky130_fd_sc_hd__xor2_1
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$7 _303_/Q _175_/Q VGND VGND VPWR VPWR final_adder.U$$7/COUT final_adder.U$$7/SUM
+ sky130_fd_sc_hd__ha_1
Xoutput302 output302/A VGND VGND VPWR VPWR o[25] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_1 U$$3383/X U$$3516/X U$$3649/X VGND VGND VPWR VPWR dadda_fa_3_93_0/CIN
+ dadda_fa_3_92_2/CIN sky130_fd_sc_hd__fa_1
Xoutput313 output313/A VGND VGND VPWR VPWR o[35] sky130_fd_sc_hd__buf_2
Xoutput324 output324/A VGND VGND VPWR VPWR o[45] sky130_fd_sc_hd__buf_2
XFILLER_126_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput335 output335/A VGND VGND VPWR VPWR o[55] sky130_fd_sc_hd__buf_2
XFILLER_160_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput346 output346/A VGND VGND VPWR VPWR o[65] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_85_0 U$$3901/X U$$4034/X U$$4167/X VGND VGND VPWR VPWR dadda_fa_3_86_0/B
+ dadda_fa_3_85_2/B sky130_fd_sc_hd__fa_1
Xoutput357 output357/A VGND VGND VPWR VPWR o[75] sky130_fd_sc_hd__buf_2
Xoutput368 output368/A VGND VGND VPWR VPWR o[85] sky130_fd_sc_hd__buf_2
Xoutput379 output379/A VGND VGND VPWR VPWR o[95] sky130_fd_sc_hd__buf_2
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_48_7 U$$2896/X U$$3029/X VGND VGND VPWR VPWR dadda_fa_2_49_3/B dadda_fa_3_48_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_141_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_61_7 dadda_fa_1_61_7/A dadda_fa_1_61_7/B dadda_fa_1_61_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_62_2/CIN dadda_fa_2_61_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_54_6 U$$3174/X U$$3307/X U$$3440/X VGND VGND VPWR VPWR dadda_fa_2_55_2/B
+ dadda_fa_2_54_5/B sky130_fd_sc_hd__fa_1
XFILLER_110_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_47_5 U$$2096/X U$$2229/X U$$2362/X VGND VGND VPWR VPWR dadda_fa_2_48_3/A
+ dadda_fa_2_47_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_6_0 dadda_fa_7_6_0/A dadda_fa_7_6_0/B dadda_fa_7_6_0/CIN VGND VGND VPWR
+ VPWR _303_/D _174_/D sky130_fd_sc_hd__fa_1
XFILLER_42_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_84_0 dadda_fa_7_84_0/A dadda_fa_7_84_0/B dadda_fa_7_84_0/CIN VGND VGND
+ VPWR VPWR _381_/D _252_/D sky130_fd_sc_hd__fa_1
XFILLER_164_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_985 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1505 input14/X VGND VGND VPWR VPWR U$$1491/B sky130_fd_sc_hd__buf_12
Xfanout1516 U$$4271/A1 VGND VGND VPWR VPWR U$$981/B1 sky130_fd_sc_hd__buf_4
Xfanout1527 U$$979/B1 VGND VGND VPWR VPWR U$$22/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout540 U$$2744/X VGND VGND VPWR VPWR U$$2844/A2 sky130_fd_sc_hd__buf_4
Xfanout1538 input125/X VGND VGND VPWR VPWR U$$3580/B1 sky130_fd_sc_hd__buf_4
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout551 U$$2679/A2 VGND VGND VPWR VPWR U$$2733/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1549 U$$4516/A1 VGND VGND VPWR VPWR U$$4377/B1 sky130_fd_sc_hd__buf_4
Xfanout562 U$$2407/A2 VGND VGND VPWR VPWR U$$2395/A2 sky130_fd_sc_hd__buf_4
XU$$4008 U$$4008/A U$$4058/B VGND VGND VPWR VPWR U$$4008/X sky130_fd_sc_hd__xor2_1
XFILLER_59_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4019 U$$4291/B1 U$$4043/A2 U$$4158/A1 U$$4043/B2 VGND VGND VPWR VPWR U$$4020/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout573 U$$2282/A2 VGND VGND VPWR VPWR U$$2248/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout584 U$$2059/X VGND VGND VPWR VPWR U$$2181/A2 sky130_fd_sc_hd__buf_6
XFILLER_76_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout595 U$$1859/A2 VGND VGND VPWR VPWR U$$1831/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3307 U$$3307/A U$$3349/B VGND VGND VPWR VPWR U$$3307/X sky130_fd_sc_hd__xor2_1
XU$$3318 U$$4001/B1 U$$3338/A2 U$$852/B1 U$$3338/B2 VGND VGND VPWR VPWR U$$3319/A
+ sky130_fd_sc_hd__a22o_1
XU$$3329 U$$3329/A U$$3335/B VGND VGND VPWR VPWR U$$3329/X sky130_fd_sc_hd__xor2_1
XFILLER_73_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2606 U$$2740/A U$$2606/B VGND VGND VPWR VPWR U$$2606/X sky130_fd_sc_hd__and2_1
XU$$2617 U$$2754/A1 U$$2665/A2 U$$2891/B1 U$$2665/B2 VGND VGND VPWR VPWR U$$2618/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2628 U$$2628/A U$$2662/B VGND VGND VPWR VPWR U$$2628/X sky130_fd_sc_hd__xor2_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2639 U$$447/A1 U$$2679/A2 U$$447/B1 U$$2679/B2 VGND VGND VPWR VPWR U$$2640/A sky130_fd_sc_hd__a22o_1
XU$$1905 U$$2042/A1 U$$1911/A2 U$$2179/B1 U$$1911/B2 VGND VGND VPWR VPWR U$$1906/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1916 U$$1916/A U$$1916/B VGND VGND VPWR VPWR U$$1916/X sky130_fd_sc_hd__xor2_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1927 U$$1927/A U$$1963/B VGND VGND VPWR VPWR U$$1927/X sky130_fd_sc_hd__xor2_1
XFILLER_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1938 U$$20/A1 U$$1980/A2 U$$22/A1 U$$1980/B2 VGND VGND VPWR VPWR U$$1939/A sky130_fd_sc_hd__a22o_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1949 U$$1949/A U$$2007/B VGND VGND VPWR VPWR U$$1949/X sky130_fd_sc_hd__xor2_1
X_404_ _405_/CLK _404_/D VGND VGND VPWR VPWR _404_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_335_ _344_/CLK _335_/D VGND VGND VPWR VPWR _335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_266_ _397_/CLK _266_/D VGND VGND VPWR VPWR _266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_197_ _344_/CLK _197_/D VGND VGND VPWR VPWR _197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_64_5 dadda_fa_2_64_5/A dadda_fa_2_64_5/B dadda_fa_2_64_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_2/A dadda_fa_4_64_0/A sky130_fd_sc_hd__fa_2
XFILLER_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_57_4 dadda_fa_2_57_4/A dadda_fa_2_57_4/B dadda_fa_2_57_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_1/CIN dadda_fa_3_57_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_49_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$12 U$$12/A1 U$$8/A2 U$$14/A1 U$$8/B2 VGND VGND VPWR VPWR U$$13/A sky130_fd_sc_hd__a22o_1
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$23 U$$23/A U$$9/B VGND VGND VPWR VPWR U$$23/X sky130_fd_sc_hd__xor2_1
XU$$34 U$$34/A1 U$$74/A2 U$$36/A1 U$$74/B2 VGND VGND VPWR VPWR U$$35/A sky130_fd_sc_hd__a22o_1
XU$$3830 U$$3830/A U$$3835/A VGND VGND VPWR VPWR U$$3830/X sky130_fd_sc_hd__xor2_1
XU$$3841 U$$3839/B U$$3836/A input52/X U$$3836/Y VGND VGND VPWR VPWR U$$3841/X sky130_fd_sc_hd__a22o_2
XU$$45 U$$45/A U$$77/B VGND VGND VPWR VPWR U$$45/X sky130_fd_sc_hd__xor2_1
XFILLER_37_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$56 U$$56/A1 U$$86/A2 U$$56/B1 U$$86/B2 VGND VGND VPWR VPWR U$$57/A sky130_fd_sc_hd__a22o_1
XU$$67 U$$67/A U$$97/B VGND VGND VPWR VPWR U$$67/X sky130_fd_sc_hd__xor2_1
XU$$3852 U$$4400/A1 U$$3892/A2 U$$4400/B1 U$$3892/B2 VGND VGND VPWR VPWR U$$3853/A
+ sky130_fd_sc_hd__a22o_1
XU$$3863 U$$3863/A U$$3867/B VGND VGND VPWR VPWR U$$3863/X sky130_fd_sc_hd__xor2_1
XFILLER_80_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$78 U$$78/A1 U$$80/A2 U$$80/A1 U$$80/B2 VGND VGND VPWR VPWR U$$79/A sky130_fd_sc_hd__a22o_1
XU$$3874 U$$4011/A1 U$$3924/A2 U$$4150/A1 U$$3924/B2 VGND VGND VPWR VPWR U$$3875/A
+ sky130_fd_sc_hd__a22o_1
XU$$89 U$$89/A U$$97/B VGND VGND VPWR VPWR U$$89/X sky130_fd_sc_hd__xor2_1
XU$$3885 U$$3885/A U$$3965/B VGND VGND VPWR VPWR U$$3885/X sky130_fd_sc_hd__xor2_1
XU$$3896 U$$4307/A1 U$$3906/A2 U$$4307/B1 U$$3906/B2 VGND VGND VPWR VPWR U$$3897/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_44_clk _218_/CLK VGND VGND VPWR VPWR _342_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_52_3 U$$1574/X U$$1707/X U$$1840/X VGND VGND VPWR VPWR dadda_fa_2_53_1/B
+ dadda_fa_2_52_4/B sky130_fd_sc_hd__fa_1
XFILLER_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_45_2 U$$895/X U$$1028/X U$$1161/X VGND VGND VPWR VPWR dadda_fa_2_46_2/CIN
+ dadda_fa_2_45_5/A sky130_fd_sc_hd__fa_1
XFILLER_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_22_1 dadda_fa_4_22_1/A dadda_fa_4_22_1/B dadda_fa_4_22_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_23_0/B dadda_fa_5_22_1/B sky130_fd_sc_hd__fa_1
XFILLER_71_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_38_1 U$$482/X U$$615/X U$$748/X VGND VGND VPWR VPWR dadda_fa_2_39_4/CIN
+ dadda_fa_2_38_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_clk _388_/CLK VGND VGND VPWR VPWR _367_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_4_15_0 U$$303/X U$$436/X U$$569/X VGND VGND VPWR VPWR dadda_fa_5_16_0/A
+ dadda_fa_5_15_1/A sky130_fd_sc_hd__fa_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1017 final_adder.U$$8/SUM final_adder.U$$503/X final_adder.U$$8/COUT
+ VGND VGND VPWR VPWR final_adder.U$$1033/B sky130_fd_sc_hd__a21o_1
XFILLER_165_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1028 final_adder.U$$4/SUM final_adder.U$$381/X VGND VGND VPWR VPWR
+ output329/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1039 final_adder.U$$240/B final_adder.U$$1039/B VGND VGND VPWR VPWR
+ output291/A sky130_fd_sc_hd__xor2_1
XFILLER_165_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1302 fanout1309/X VGND VGND VPWR VPWR U$$3907/B sky130_fd_sc_hd__buf_6
XFILLER_121_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_67_3 dadda_fa_3_67_3/A dadda_fa_3_67_3/B dadda_fa_3_67_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_1/B dadda_fa_4_67_2/CIN sky130_fd_sc_hd__fa_1
Xfanout1313 U$$3792/B VGND VGND VPWR VPWR U$$3740/B sky130_fd_sc_hd__buf_6
XFILLER_79_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1324 U$$907/B VGND VGND VPWR VPWR U$$913/B sky130_fd_sc_hd__buf_4
Xfanout1335 U$$3659/B VGND VGND VPWR VPWR U$$3698/A sky130_fd_sc_hd__buf_4
XFILLER_120_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1346 input44/X VGND VGND VPWR VPWR U$$3335/B sky130_fd_sc_hd__buf_6
Xfanout1357 fanout1364/X VGND VGND VPWR VPWR U$$3242/B sky130_fd_sc_hd__buf_6
Xfanout1368 input40/X VGND VGND VPWR VPWR U$$3151/A sky130_fd_sc_hd__buf_4
Xfanout1379 U$$2986/B VGND VGND VPWR VPWR U$$3004/B sky130_fd_sc_hd__buf_6
Xfanout392 U$$902/A2 VGND VGND VPWR VPWR U$$898/A2 sky130_fd_sc_hd__buf_4
XFILLER_87_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3104 U$$3239/B1 U$$3108/A2 U$$3106/A1 U$$3108/B2 VGND VGND VPWR VPWR U$$3105/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3115 U$$3115/A U$$3119/B VGND VGND VPWR VPWR U$$3115/X sky130_fd_sc_hd__xor2_1
XU$$3126 U$$3948/A1 U$$3148/A2 U$$251/A1 U$$3148/B2 VGND VGND VPWR VPWR U$$3127/A
+ sky130_fd_sc_hd__a22o_1
XU$$3137 U$$3137/A U$$3147/B VGND VGND VPWR VPWR U$$3137/X sky130_fd_sc_hd__xor2_1
XU$$2403 U$$620/B1 U$$2407/A2 U$$487/A1 U$$2407/B2 VGND VGND VPWR VPWR U$$2404/A sky130_fd_sc_hd__a22o_1
XU$$3148 U$$3285/A1 U$$3148/A2 U$$3148/B1 U$$3148/B2 VGND VGND VPWR VPWR U$$3149/A
+ sky130_fd_sc_hd__a22o_1
XU$$3159 U$$4392/A1 U$$3199/A2 U$$3296/B1 U$$3199/B2 VGND VGND VPWR VPWR U$$3160/A
+ sky130_fd_sc_hd__a22o_1
XU$$2414 U$$2414/A U$$2416/B VGND VGND VPWR VPWR U$$2414/X sky130_fd_sc_hd__xor2_1
XU$$2425 U$$3110/A1 U$$2445/A2 U$$3112/A1 U$$2445/B2 VGND VGND VPWR VPWR U$$2426/A
+ sky130_fd_sc_hd__a22o_1
XU$$2436 U$$2436/A U$$2466/A VGND VGND VPWR VPWR U$$2436/X sky130_fd_sc_hd__xor2_1
XU$$1702 U$$880/A1 U$$1702/A2 U$$882/A1 U$$1702/B2 VGND VGND VPWR VPWR U$$1703/A sky130_fd_sc_hd__a22o_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2447 U$$4365/A1 U$$2459/A2 U$$4365/B1 U$$2459/B2 VGND VGND VPWR VPWR U$$2448/A
+ sky130_fd_sc_hd__a22o_1
XU$$1713 U$$1713/A U$$1721/B VGND VGND VPWR VPWR U$$1713/X sky130_fd_sc_hd__xor2_1
XU$$2458 U$$2458/A U$$2465/A VGND VGND VPWR VPWR U$$2458/X sky130_fd_sc_hd__xor2_1
XU$$2469 U$$2575/B U$$2469/B VGND VGND VPWR VPWR U$$2469/X sky130_fd_sc_hd__and2_1
XU$$1724 U$$902/A1 U$$1726/A2 U$$765/B1 U$$1726/B2 VGND VGND VPWR VPWR U$$1725/A sky130_fd_sc_hd__a22o_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1735 U$$1735/A U$$1741/B VGND VGND VPWR VPWR U$$1735/X sky130_fd_sc_hd__xor2_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1746 U$$787/A1 U$$1758/A2 U$$787/B1 U$$1758/B2 VGND VGND VPWR VPWR U$$1747/A sky130_fd_sc_hd__a22o_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$408_1830 VGND VGND VPWR VPWR U$$408_1830/HI U$$408/B1 sky130_fd_sc_hd__conb_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1757 U$$1757/A U$$1761/B VGND VGND VPWR VPWR U$$1757/X sky130_fd_sc_hd__xor2_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1768 U$$2042/A1 U$$1774/A2 U$$2179/B1 U$$1774/B2 VGND VGND VPWR VPWR U$$1769/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1779 U$$1779/A U$$1781/A VGND VGND VPWR VPWR U$$1779/X sky130_fd_sc_hd__xor2_1
XFILLER_42_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_318_ _321_/CLK _318_/D VGND VGND VPWR VPWR _318_/Q sky130_fd_sc_hd__dfxtp_1
Xinput12 a[1] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__buf_4
Xinput23 a[2] VGND VGND VPWR VPWR U$$138/A sky130_fd_sc_hd__buf_2
XFILLER_174_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput34 a[3] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__buf_4
Xinput45 a[4] VGND VGND VPWR VPWR U$$275/A sky130_fd_sc_hd__buf_2
X_249_ _382_/CLK _249_/D VGND VGND VPWR VPWR _249_/Q sky130_fd_sc_hd__dfxtp_1
Xinput56 a[5] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__buf_6
XFILLER_155_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput67 b[11] VGND VGND VPWR VPWR input67/X sky130_fd_sc_hd__buf_2
Xinput78 b[21] VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput89 b[31] VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_62_2 dadda_fa_2_62_2/A dadda_fa_2_62_2/B dadda_fa_2_62_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_1/A dadda_fa_3_62_3/A sky130_fd_sc_hd__fa_1
XFILLER_69_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$409 final_adder.U$$408/B final_adder.U$$287/X final_adder.U$$283/X
+ VGND VGND VPWR VPWR final_adder.U$$409/X sky130_fd_sc_hd__a21o_1
XFILLER_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_55_1 dadda_fa_2_55_1/A dadda_fa_2_55_1/B dadda_fa_2_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_0/CIN dadda_fa_3_55_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_32_0 dadda_fa_5_32_0/A dadda_fa_5_32_0/B dadda_fa_5_32_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_33_0/A dadda_fa_6_32_0/CIN sky130_fd_sc_hd__fa_1
XU$$4350 U$$4350/A U$$4350/B VGND VGND VPWR VPWR U$$4350/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_48_0 U$$3162/X U$$3295/X U$$3335/B VGND VGND VPWR VPWR dadda_fa_3_49_0/B
+ dadda_fa_3_48_2/B sky130_fd_sc_hd__fa_1
XU$$4361 U$$4361/A1 U$$4369/A2 U$$4363/A1 U$$4369/B2 VGND VGND VPWR VPWR U$$4362/A
+ sky130_fd_sc_hd__a22o_1
XU$$4372 U$$4372/A U$$4374/B VGND VGND VPWR VPWR U$$4372/X sky130_fd_sc_hd__xor2_1
XU$$4383 U$$4383/A VGND VGND VPWR VPWR U$$4383/Y sky130_fd_sc_hd__inv_1
XU$$4394 input76/X U$$4388/X U$$4396/A1 U$$4428/B2 VGND VGND VPWR VPWR U$$4395/A sky130_fd_sc_hd__a22o_1
XU$$3660 U$$4345/A1 U$$3682/A2 U$$4482/B1 U$$3682/B2 VGND VGND VPWR VPWR U$$3661/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3671 U$$3671/A U$$3681/B VGND VGND VPWR VPWR U$$3671/X sky130_fd_sc_hd__xor2_1
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3682 U$$3817/B1 U$$3682/A2 U$$3684/A1 U$$3682/B2 VGND VGND VPWR VPWR U$$3683/A
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_17_clk _370_/CLK VGND VGND VPWR VPWR _402_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3693 U$$3693/A U$$3698/A VGND VGND VPWR VPWR U$$3693/X sky130_fd_sc_hd__xor2_1
XFILLER_34_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2970 U$$2970/A U$$2974/B VGND VGND VPWR VPWR U$$2970/X sky130_fd_sc_hd__xor2_1
XU$$2981 U$$4486/B1 U$$3011/A2 U$$4353/A1 U$$3011/B2 VGND VGND VPWR VPWR U$$2982/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_9_1 input256/X dadda_fa_5_9_1/B dadda_ha_4_9_0/SUM VGND VGND VPWR VPWR
+ dadda_fa_6_10_0/B dadda_fa_7_9_0/A sky130_fd_sc_hd__fa_1
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2992 U$$2992/A U$$3004/B VGND VGND VPWR VPWR U$$2992/X sky130_fd_sc_hd__xor2_1
XFILLER_33_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_77_2 dadda_fa_4_77_2/A dadda_fa_4_77_2/B dadda_fa_4_77_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_78_0/CIN dadda_fa_5_77_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_47_0 dadda_fa_7_47_0/A dadda_fa_7_47_0/B dadda_fa_7_47_0/CIN VGND VGND
+ VPWR VPWR _344_/D _215_/D sky130_fd_sc_hd__fa_2
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$921 final_adder.U$$150/A final_adder.U$$859/X final_adder.U$$921/B1
+ VGND VGND VPWR VPWR final_adder.U$$921/X sky130_fd_sc_hd__a21o_1
XFILLER_69_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$943 final_adder.U$$172/A final_adder.U$$881/X final_adder.U$$943/B1
+ VGND VGND VPWR VPWR final_adder.U$$943/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_0 U$$107/X U$$240/X U$$373/X VGND VGND VPWR VPWR dadda_fa_2_51_0/B
+ dadda_fa_2_50_3/B sky130_fd_sc_hd__fa_1
XFILLER_113_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$965 final_adder.U$$194/A final_adder.U$$807/X final_adder.U$$965/B1
+ VGND VGND VPWR VPWR final_adder.U$$965/X sky130_fd_sc_hd__a21o_1
XU$$804 U$$804/A U$$804/B VGND VGND VPWR VPWR U$$804/X sky130_fd_sc_hd__xor2_1
XU$$815 U$$952/A1 U$$817/A2 U$$954/A1 U$$817/B2 VGND VGND VPWR VPWR U$$816/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$987 final_adder.U$$216/A final_adder.U$$829/X final_adder.U$$987/B1
+ VGND VGND VPWR VPWR final_adder.U$$987/X sky130_fd_sc_hd__a21o_1
XU$$826 U$$824/Y input4/X U$$822/A U$$825/X U$$822/Y VGND VGND VPWR VPWR U$$826/X
+ sky130_fd_sc_hd__a32o_1
XU$$837 U$$837/A U$$907/B VGND VGND VPWR VPWR U$$837/X sky130_fd_sc_hd__xor2_1
XU$$848 U$$985/A1 U$$904/A2 U$$987/A1 U$$904/B2 VGND VGND VPWR VPWR U$$849/A sky130_fd_sc_hd__a22o_1
XU$$859 U$$859/A U$$895/B VGND VGND VPWR VPWR U$$859/X sky130_fd_sc_hd__xor2_1
XU$$1009 U$$50/A1 U$$979/A2 U$$50/B1 U$$979/B2 VGND VGND VPWR VPWR U$$1010/A sky130_fd_sc_hd__a22o_1
XFILLER_106_1003 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_72_1 dadda_fa_3_72_1/A dadda_fa_3_72_1/B dadda_fa_3_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_0/CIN dadda_fa_4_72_2/A sky130_fd_sc_hd__fa_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1110 U$$52/A1 VGND VGND VPWR VPWR U$$598/B1 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_3_65_0 dadda_fa_3_65_0/A dadda_fa_3_65_0/B dadda_fa_3_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_0/B dadda_fa_4_65_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_26_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1121 U$$872/A1 VGND VGND VPWR VPWR U$$50/A1 sky130_fd_sc_hd__buf_4
XFILLER_39_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1132 U$$3884/A1 VGND VGND VPWR VPWR U$$4432/A1 sky130_fd_sc_hd__buf_6
XFILLER_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1143 U$$2923/A1 VGND VGND VPWR VPWR U$$868/A1 sky130_fd_sc_hd__buf_4
XFILLER_121_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1154 input74/X VGND VGND VPWR VPWR U$$4291/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1165 U$$4152/A1 VGND VGND VPWR VPWR U$$40/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1176 input72/X VGND VGND VPWR VPWR U$$4424/A1 sky130_fd_sc_hd__buf_4
Xfanout1187 U$$3870/B1 VGND VGND VPWR VPWR U$$721/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1198 U$$982/B VGND VGND VPWR VPWR U$$1046/B sky130_fd_sc_hd__clkbuf_4
XFILLER_75_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2200 U$$967/A1 U$$2252/A2 U$$969/A1 U$$2252/B2 VGND VGND VPWR VPWR U$$2201/A sky130_fd_sc_hd__a22o_1
XFILLER_47_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2211 U$$2211/A U$$2253/B VGND VGND VPWR VPWR U$$2211/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_101_1 dadda_fa_4_101_1/A dadda_fa_4_101_1/B dadda_fa_4_101_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_102_0/B dadda_fa_5_101_1/B sky130_fd_sc_hd__fa_1
XU$$2222 U$$989/A1 U$$2254/A2 U$$991/A1 U$$2254/B2 VGND VGND VPWR VPWR U$$2223/A sky130_fd_sc_hd__a22o_1
XFILLER_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2233 U$$2233/A U$$2269/B VGND VGND VPWR VPWR U$$2233/X sky130_fd_sc_hd__xor2_1
XU$$2244 U$$874/A1 U$$2282/A2 U$$876/A1 U$$2282/B2 VGND VGND VPWR VPWR U$$2245/A sky130_fd_sc_hd__a22o_1
XU$$1510 U$$1644/A U$$1510/B VGND VGND VPWR VPWR U$$1510/X sky130_fd_sc_hd__and2_1
XU$$2255 U$$2255/A U$$2269/B VGND VGND VPWR VPWR U$$2255/X sky130_fd_sc_hd__xor2_1
XFILLER_90_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1521 U$$2754/A1 U$$1563/A2 U$$2891/B1 U$$1563/B2 VGND VGND VPWR VPWR U$$1522/A
+ sky130_fd_sc_hd__a22o_1
XU$$2266 U$$3499/A1 U$$2310/A2 U$$3775/A1 U$$2310/B2 VGND VGND VPWR VPWR U$$2267/A
+ sky130_fd_sc_hd__a22o_1
XU$$1532 U$$1532/A U$$1568/B VGND VGND VPWR VPWR U$$1532/X sky130_fd_sc_hd__xor2_1
XU$$2277 U$$2277/A U$$2327/B VGND VGND VPWR VPWR U$$2277/X sky130_fd_sc_hd__xor2_1
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1543 U$$36/A1 U$$1575/A2 U$$38/A1 U$$1575/B2 VGND VGND VPWR VPWR U$$1544/A sky130_fd_sc_hd__a22o_1
XU$$2288 U$$4478/B1 U$$2326/A2 U$$4345/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2289/A
+ sky130_fd_sc_hd__a22o_1
XU$$1554 U$$1554/A U$$1564/B VGND VGND VPWR VPWR U$$1554/X sky130_fd_sc_hd__xor2_1
XU$$2299 U$$2299/A U$$2301/B VGND VGND VPWR VPWR U$$2299/X sky130_fd_sc_hd__xor2_1
XU$$1565 U$$56/B1 U$$1567/A2 U$$469/B1 U$$1567/B2 VGND VGND VPWR VPWR U$$1566/A sky130_fd_sc_hd__a22o_1
XU$$1576 U$$1576/A U$$1584/B VGND VGND VPWR VPWR U$$1576/X sky130_fd_sc_hd__xor2_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1587 U$$900/B1 U$$1587/A2 U$$765/B1 U$$1587/B2 VGND VGND VPWR VPWR U$$1588/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_7_122_0 dadda_fa_7_122_0/A dadda_fa_7_122_0/B dadda_fa_7_122_0/CIN VGND
+ VGND VPWR VPWR _419_/D _290_/D sky130_fd_sc_hd__fa_1
XU$$1598 U$$1598/A U$$1608/B VGND VGND VPWR VPWR U$$1598/X sky130_fd_sc_hd__xor2_1
XFILLER_42_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_87_1 dadda_fa_5_87_1/A dadda_fa_5_87_1/B dadda_fa_5_87_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_88_0/B dadda_fa_7_87_0/A sky130_fd_sc_hd__fa_2
XFILLER_131_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4511_1903 VGND VGND VPWR VPWR U$$4511_1903/HI U$$4511/B sky130_fd_sc_hd__conb_1
XFILLER_131_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_79_8 U$$4288/X U$$4421/X input233/X VGND VGND VPWR VPWR dadda_fa_2_80_3/A
+ dadda_fa_3_79_0/A sky130_fd_sc_hd__fa_2
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$206 final_adder.U$$206/A final_adder.U$$206/B VGND VGND VPWR VPWR
+ final_adder.U$$334/B sky130_fd_sc_hd__and2_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$217 final_adder.U$$216/B final_adder.U$$987/B1 final_adder.U$$217/B1
+ VGND VGND VPWR VPWR final_adder.U$$217/X sky130_fd_sc_hd__a21o_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$228 final_adder.U$$228/A final_adder.U$$228/B VGND VGND VPWR VPWR
+ final_adder.U$$356/B sky130_fd_sc_hd__and2_1
XFILLER_100_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$239 final_adder.U$$238/B final_adder.U$$239/A2 final_adder.U$$239/B1
+ VGND VGND VPWR VPWR final_adder.U$$239/X sky130_fd_sc_hd__a21o_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4180 U$$4454/A1 U$$4240/A2 U$$4456/A1 U$$4240/B2 VGND VGND VPWR VPWR U$$4181/A
+ sky130_fd_sc_hd__a22o_1
XU$$4191 U$$4191/A U$$4191/B VGND VGND VPWR VPWR U$$4191/X sky130_fd_sc_hd__xor2_1
XU$$3490 U$$3490/A U$$3506/B VGND VGND VPWR VPWR U$$3490/X sky130_fd_sc_hd__xor2_1
XFILLER_129_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_82_0 dadda_fa_4_82_0/A dadda_fa_4_82_0/B dadda_fa_4_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_83_0/A dadda_fa_5_82_1/A sky130_fd_sc_hd__fa_1
XFILLER_146_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_103_3 dadda_fa_3_103_3/A dadda_fa_3_103_3/B dadda_fa_3_103_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_104_1/B dadda_fa_4_103_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_150_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput202 c[50] VGND VGND VPWR VPWR input202/X sky130_fd_sc_hd__clkbuf_2
Xinput213 c[60] VGND VGND VPWR VPWR input213/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput224 c[70] VGND VGND VPWR VPWR input224/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput235 c[80] VGND VGND VPWR VPWR input235/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput246 c[90] VGND VGND VPWR VPWR input246/X sky130_fd_sc_hd__buf_2
XFILLER_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$740 final_adder.U$$772/B final_adder.U$$740/B VGND VGND VPWR VPWR
+ final_adder.U$$740/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$751 final_adder.U$$750/B final_adder.U$$671/X final_adder.U$$639/X
+ VGND VGND VPWR VPWR final_adder.U$$751/X sky130_fd_sc_hd__a21o_1
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$762 final_adder.U$$794/B final_adder.U$$762/B VGND VGND VPWR VPWR
+ final_adder.U$$762/X sky130_fd_sc_hd__and2_1
XU$$601 U$$601/A U$$637/B VGND VGND VPWR VPWR U$$601/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$773 final_adder.U$$772/B final_adder.U$$693/X final_adder.U$$661/X
+ VGND VGND VPWR VPWR final_adder.U$$773/X sky130_fd_sc_hd__a21o_1
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$612 U$$612/A1 U$$642/A2 U$$612/B1 U$$642/B2 VGND VGND VPWR VPWR U$$613/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$784 final_adder.U$$784/A final_adder.U$$784/B VGND VGND VPWR VPWR
+ final_adder.U$$784/X sky130_fd_sc_hd__and2_1
XFILLER_17_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$623 U$$623/A U$$631/B VGND VGND VPWR VPWR U$$623/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$795 final_adder.U$$794/B final_adder.U$$715/X final_adder.U$$683/X
+ VGND VGND VPWR VPWR final_adder.U$$795/X sky130_fd_sc_hd__a21o_1
XU$$634 U$$86/A1 U$$636/A2 U$$88/A1 U$$636/B2 VGND VGND VPWR VPWR U$$635/A sky130_fd_sc_hd__a22o_1
XFILLER_84_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$645 U$$645/A U$$684/A VGND VGND VPWR VPWR U$$645/X sky130_fd_sc_hd__xor2_1
XU$$656 U$$930/A1 U$$674/A2 U$$932/A1 U$$674/B2 VGND VGND VPWR VPWR U$$657/A sky130_fd_sc_hd__a22o_1
XU$$667 U$$667/A U$$669/B VGND VGND VPWR VPWR U$$667/X sky130_fd_sc_hd__xor2_1
XU$$678 U$$678/A1 U$$682/A2 U$$678/B1 U$$682/B2 VGND VGND VPWR VPWR U$$679/A sky130_fd_sc_hd__a22o_1
XU$$689 U$$687/Y input2/X U$$685/A U$$688/X U$$685/Y VGND VGND VPWR VPWR U$$689/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_72_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_97_0 dadda_fa_6_97_0/A dadda_fa_6_97_0/B dadda_fa_6_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_98_0/B dadda_fa_7_97_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_2_33_5 U$$2068/X U$$2201/X VGND VGND VPWR VPWR dadda_fa_3_34_2/A dadda_fa_4_33_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_67_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_32_3 U$$1268/X U$$1401/X U$$1534/X VGND VGND VPWR VPWR dadda_fa_3_33_1/B
+ dadda_fa_3_32_3/B sky130_fd_sc_hd__fa_1
XU$$2030 U$$2576/B1 U$$2046/A2 U$$936/A1 U$$2046/B2 VGND VGND VPWR VPWR U$$2031/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2041 U$$2041/A U$$2043/B VGND VGND VPWR VPWR U$$2041/X sky130_fd_sc_hd__xor2_1
XFILLER_90_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2052 U$$3833/A1 U$$2052/A2 U$$2052/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2053/A
+ sky130_fd_sc_hd__a22o_1
XU$$2063 U$$3022/A1 U$$2139/A2 U$$3022/B1 U$$2139/B2 VGND VGND VPWR VPWR U$$2064/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2074 U$$2074/A U$$2106/B VGND VGND VPWR VPWR U$$2074/X sky130_fd_sc_hd__xor2_1
XU$$1340 U$$1340/A U$$1364/B VGND VGND VPWR VPWR U$$1340/X sky130_fd_sc_hd__xor2_1
XU$$2085 U$$989/A1 U$$2097/A2 U$$989/B1 U$$2097/B2 VGND VGND VPWR VPWR U$$2086/A sky130_fd_sc_hd__a22o_1
XU$$2096 U$$2096/A U$$2096/B VGND VGND VPWR VPWR U$$2096/X sky130_fd_sc_hd__xor2_1
XU$$1351 U$$253/B1 U$$1353/A2 U$$120/A1 U$$1353/B2 VGND VGND VPWR VPWR U$$1352/A sky130_fd_sc_hd__a22o_1
XU$$1362 U$$1362/A U$$1364/B VGND VGND VPWR VPWR U$$1362/X sky130_fd_sc_hd__xor2_1
XU$$1373 U$$1507/A U$$1373/B VGND VGND VPWR VPWR U$$1373/X sky130_fd_sc_hd__and2_1
XU$$1384 U$$2480/A1 U$$1432/A2 U$$3030/A1 U$$1432/B2 VGND VGND VPWR VPWR U$$1385/A
+ sky130_fd_sc_hd__a22o_1
XU$$1395 U$$1395/A U$$1427/B VGND VGND VPWR VPWR U$$1395/X sky130_fd_sc_hd__xor2_1
XFILLER_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout903 U$$1238/X VGND VGND VPWR VPWR U$$1353/B2 sky130_fd_sc_hd__buf_6
XFILLER_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout914 U$$102/B2 VGND VGND VPWR VPWR U$$98/B2 sky130_fd_sc_hd__buf_4
Xfanout925 U$$4502/B2 VGND VGND VPWR VPWR U$$4506/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_77_5 U$$3353/X U$$3486/X U$$3619/X VGND VGND VPWR VPWR dadda_fa_2_78_2/A
+ dadda_fa_2_77_5/A sky130_fd_sc_hd__fa_1
Xfanout936 U$$910/A1 VGND VGND VPWR VPWR U$$3650/A1 sky130_fd_sc_hd__buf_6
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout947 U$$4398/A1 VGND VGND VPWR VPWR U$$3713/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout958 fanout966/X VGND VGND VPWR VPWR U$$632/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_58_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout969 U$$3642/B1 VGND VGND VPWR VPWR U$$3370/A1 sky130_fd_sc_hd__buf_4
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$80 _376_/Q _248_/Q VGND VGND VPWR VPWR final_adder.U$$945/B1 final_adder.U$$174/A
+ sky130_fd_sc_hd__ha_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$91 _387_/Q _259_/Q VGND VGND VPWR VPWR final_adder.U$$165/B1 final_adder.U$$164/B
+ sky130_fd_sc_hd__ha_1
XFILLER_110_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_86_0_1926 VGND VGND VPWR VPWR dadda_fa_1_86_0/A dadda_fa_1_86_0_1926/LO
+ sky130_fd_sc_hd__conb_1
Xdadda_fa_3_101_0 U$$4199/X U$$4332/X U$$4465/X VGND VGND VPWR VPWR dadda_fa_4_102_0/B
+ dadda_fa_4_101_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_65_3 U$$1334/X U$$1467/X U$$1600/X VGND VGND VPWR VPWR dadda_fa_1_66_6/B
+ dadda_fa_1_65_8/B sky130_fd_sc_hd__fa_1
XFILLER_77_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_42_2 dadda_fa_3_42_2/A dadda_fa_3_42_2/B dadda_fa_3_42_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_1/A dadda_fa_4_42_2/B sky130_fd_sc_hd__fa_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_58_2 U$$921/X U$$1054/X U$$1187/X VGND VGND VPWR VPWR dadda_fa_1_59_7/B
+ dadda_fa_1_58_8/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$570 final_adder.U$$578/B final_adder.U$$570/B VGND VGND VPWR VPWR
+ final_adder.U$$690/B sky130_fd_sc_hd__and2_1
Xdadda_fa_3_35_1 dadda_fa_3_35_1/A dadda_fa_3_35_1/B dadda_fa_3_35_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_0/CIN dadda_fa_4_35_2/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$581 final_adder.U$$580/B final_adder.U$$465/X final_adder.U$$457/X
+ VGND VGND VPWR VPWR final_adder.U$$581/X sky130_fd_sc_hd__a21o_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$420 U$$420/A U$$448/B VGND VGND VPWR VPWR U$$420/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$592 final_adder.U$$600/B final_adder.U$$592/B VGND VGND VPWR VPWR
+ final_adder.U$$712/B sky130_fd_sc_hd__and2_1
XU$$431 U$$20/A1 U$$447/A2 U$$22/A1 U$$447/B2 VGND VGND VPWR VPWR U$$432/A sky130_fd_sc_hd__a22o_1
XU$$442 U$$442/A U$$506/B VGND VGND VPWR VPWR U$$442/X sky130_fd_sc_hd__xor2_1
XU$$453 U$$999/B1 U$$501/A2 U$$866/A1 U$$501/B2 VGND VGND VPWR VPWR U$$454/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_12_0 dadda_fa_6_12_0/A dadda_fa_6_12_0/B dadda_fa_6_12_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_13_0/B dadda_fa_7_12_0/CIN sky130_fd_sc_hd__fa_1
XU$$464 U$$464/A U$$498/B VGND VGND VPWR VPWR U$$464/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_28_0 U$$1526/X U$$1659/X U$$1792/X VGND VGND VPWR VPWR dadda_fa_4_29_0/B
+ dadda_fa_4_28_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_45_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$475 U$$747/B1 U$$479/A2 U$$749/B1 U$$479/B2 VGND VGND VPWR VPWR U$$476/A sky130_fd_sc_hd__a22o_1
XFILLER_44_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$486 U$$486/A U$$504/B VGND VGND VPWR VPWR U$$486/X sky130_fd_sc_hd__xor2_1
XU$$497 U$$632/B1 U$$497/A2 U$$499/A1 U$$497/B2 VGND VGND VPWR VPWR U$$498/A sky130_fd_sc_hd__a22o_1
XFILLER_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_94_5 dadda_fa_2_94_5/A dadda_fa_2_94_5/B dadda_fa_2_94_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_95_2/A dadda_fa_4_94_0/A sky130_fd_sc_hd__fa_2
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_87_4 dadda_fa_2_87_4/A dadda_fa_2_87_4/B dadda_fa_2_87_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_88_1/CIN dadda_fa_3_87_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_2_24_1 U$$454/X U$$587/X VGND VGND VPWR VPWR dadda_fa_3_25_3/B dadda_fa_4_24_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_68_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_30_0 U$$67/X U$$200/X U$$333/X VGND VGND VPWR VPWR dadda_fa_3_31_1/A dadda_fa_3_30_2/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_35_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_103_2 U$$3538/X U$$3671/X U$$3804/X VGND VGND VPWR VPWR dadda_fa_3_104_3/A
+ dadda_fa_4_103_0/A sky130_fd_sc_hd__fa_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1170 U$$74/A1 U$$1170/A2 U$$74/B1 U$$1170/B2 VGND VGND VPWR VPWR U$$1171/A sky130_fd_sc_hd__a22o_1
XU$$1181 U$$1181/A U$$1227/B VGND VGND VPWR VPWR U$$1181/X sky130_fd_sc_hd__xor2_1
XU$$1192 U$$96/A1 U$$1230/A2 U$$98/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1193/A sky130_fd_sc_hd__a22o_1
XFILLER_148_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_117_0 dadda_fa_5_117_0/A dadda_fa_5_117_0/B dadda_fa_5_117_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_118_0/A dadda_fa_6_117_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_74_0_1921 VGND VGND VPWR VPWR dadda_fa_0_74_0/A dadda_fa_0_74_0_1921/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_117_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1004 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_82_3 U$$2432/X U$$2565/X U$$2698/X VGND VGND VPWR VPWR dadda_fa_2_83_2/B
+ dadda_fa_2_82_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout700 U$$416/X VGND VGND VPWR VPWR U$$545/B2 sky130_fd_sc_hd__buf_6
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout711 U$$4043/B2 VGND VGND VPWR VPWR U$$4045/B2 sky130_fd_sc_hd__buf_4
Xfanout1709 input108/X VGND VGND VPWR VPWR U$$2844/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout722 U$$3966/B2 VGND VGND VPWR VPWR U$$3970/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_75_2 U$$2418/X U$$2551/X U$$2684/X VGND VGND VPWR VPWR dadda_fa_2_76_1/A
+ dadda_fa_2_75_4/A sky130_fd_sc_hd__fa_1
XFILLER_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout733 U$$3833/B2 VGND VGND VPWR VPWR U$$3825/B2 sky130_fd_sc_hd__buf_4
Xfanout744 U$$3511/B2 VGND VGND VPWR VPWR U$$3505/B2 sky130_fd_sc_hd__buf_4
Xfanout755 U$$3293/X VGND VGND VPWR VPWR U$$3378/B2 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_4_52_1 dadda_fa_4_52_1/A dadda_fa_4_52_1/B dadda_fa_4_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_53_0/B dadda_fa_5_52_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_68_1 U$$2936/X U$$3069/X U$$3202/X VGND VGND VPWR VPWR dadda_fa_2_69_0/CIN
+ dadda_fa_2_68_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout766 U$$3251/B2 VGND VGND VPWR VPWR U$$3283/B2 sky130_fd_sc_hd__buf_4
Xfanout777 U$$3118/B2 VGND VGND VPWR VPWR U$$3144/B2 sky130_fd_sc_hd__buf_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout788 U$$279/X VGND VGND VPWR VPWR U$$352/B2 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_4_45_0 dadda_fa_4_45_0/A dadda_fa_4_45_0/B dadda_fa_4_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_46_0/A dadda_fa_5_45_1/A sky130_fd_sc_hd__fa_1
Xfanout799 U$$2745/X VGND VGND VPWR VPWR U$$2844/B2 sky130_fd_sc_hd__buf_4
XFILLER_46_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_420_ _420_/CLK _420_/D VGND VGND VPWR VPWR _420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_351_ _353_/CLK _351_/D VGND VGND VPWR VPWR _351_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_282_ _416_/CLK _282_/D VGND VGND VPWR VPWR _282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_97_3 dadda_fa_3_97_3/A dadda_fa_3_97_3/B dadda_fa_3_97_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_1/B dadda_fa_4_97_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_154_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_70_1 U$$812/X U$$945/X U$$1078/X VGND VGND VPWR VPWR dadda_fa_1_71_6/CIN
+ dadda_fa_1_70_8/A sky130_fd_sc_hd__fa_1
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_63_0 U$$133/X U$$266/X U$$399/X VGND VGND VPWR VPWR dadda_fa_1_64_5/B
+ dadda_fa_1_63_7/B sky130_fd_sc_hd__fa_1
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$250 U$$250/A U$$254/B VGND VGND VPWR VPWR U$$250/X sky130_fd_sc_hd__xor2_1
XU$$261 U$$672/A1 U$$271/A2 U$$672/B1 U$$271/B2 VGND VGND VPWR VPWR U$$262/A sky130_fd_sc_hd__a22o_1
XU$$272 U$$272/A U$$274/A VGND VGND VPWR VPWR U$$272/X sky130_fd_sc_hd__xor2_1
XFILLER_17_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$283 U$$283/A U$$313/B VGND VGND VPWR VPWR U$$283/X sky130_fd_sc_hd__xor2_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$294 U$$979/A1 U$$346/A2 U$$979/B1 U$$346/B2 VGND VGND VPWR VPWR U$$295/A sky130_fd_sc_hd__a22o_1
XFILLER_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$0 U$$0/A VGND VGND VPWR VPWR U$$0/Y sky130_fd_sc_hd__inv_1
XFILLER_118_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$8 _304_/Q _176_/Q VGND VGND VPWR VPWR final_adder.U$$8/COUT final_adder.U$$8/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_146_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput303 output303/A VGND VGND VPWR VPWR o[26] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_2 U$$3782/X U$$3915/X U$$4048/X VGND VGND VPWR VPWR dadda_fa_3_93_1/A
+ dadda_fa_3_92_3/A sky130_fd_sc_hd__fa_1
Xoutput314 output314/A VGND VGND VPWR VPWR o[36] sky130_fd_sc_hd__buf_2
XFILLER_142_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput325 output325/A VGND VGND VPWR VPWR o[46] sky130_fd_sc_hd__buf_2
Xoutput336 output336/A VGND VGND VPWR VPWR o[56] sky130_fd_sc_hd__buf_2
Xoutput347 output347/A VGND VGND VPWR VPWR o[66] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_85_1 U$$4300/X U$$4433/X input240/X VGND VGND VPWR VPWR dadda_fa_3_86_0/CIN
+ dadda_fa_3_85_2/CIN sky130_fd_sc_hd__fa_1
Xoutput358 output358/A VGND VGND VPWR VPWR o[76] sky130_fd_sc_hd__buf_2
XFILLER_160_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput369 output369/A VGND VGND VPWR VPWR o[86] sky130_fd_sc_hd__buf_2
XFILLER_99_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_62_0 dadda_fa_5_62_0/A dadda_fa_5_62_0/B dadda_fa_5_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_63_0/A dadda_fa_6_62_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_102_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_78_0 dadda_fa_2_78_0/A dadda_fa_2_78_0/B dadda_fa_2_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_0/B dadda_fa_3_78_2/B sky130_fd_sc_hd__fa_1
XFILLER_102_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_61_8 dadda_fa_1_61_8/A dadda_fa_1_61_8/B dadda_fa_1_61_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_62_3/A dadda_fa_3_61_0/A sky130_fd_sc_hd__fa_2
XFILLER_95_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_54_7 U$$3573/X U$$3706/X U$$3792/B VGND VGND VPWR VPWR dadda_fa_2_55_2/CIN
+ dadda_fa_2_54_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_77_0 dadda_fa_7_77_0/A dadda_fa_7_77_0/B dadda_fa_7_77_0/CIN VGND VGND
+ VPWR VPWR _374_/D _245_/D sky130_fd_sc_hd__fa_1
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_80_0 dadda_fa_1_80_0/A U$$1231/X U$$1364/X VGND VGND VPWR VPWR dadda_fa_2_81_0/CIN
+ dadda_fa_2_80_3/B sky130_fd_sc_hd__fa_1
Xfanout1506 U$$2629/A1 VGND VGND VPWR VPWR U$$983/B1 sky130_fd_sc_hd__buf_4
XFILLER_104_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1517 U$$4271/A1 VGND VGND VPWR VPWR U$$4132/B1 sky130_fd_sc_hd__buf_4
Xfanout530 U$$408/A2 VGND VGND VPWR VPWR U$$406/A2 sky130_fd_sc_hd__buf_4
Xfanout1528 U$$4406/A1 VGND VGND VPWR VPWR U$$979/B1 sky130_fd_sc_hd__buf_4
Xfanout1539 U$$545/A1 VGND VGND VPWR VPWR U$$406/B1 sky130_fd_sc_hd__buf_4
Xfanout541 U$$2812/A2 VGND VGND VPWR VPWR U$$2856/A2 sky130_fd_sc_hd__buf_6
Xfanout552 U$$2607/X VGND VGND VPWR VPWR U$$2679/A2 sky130_fd_sc_hd__buf_4
Xfanout563 U$$2445/A2 VGND VGND VPWR VPWR U$$2407/A2 sky130_fd_sc_hd__buf_6
XU$$4009 U$$4283/A1 U$$4057/A2 U$$4011/A1 U$$4057/B2 VGND VGND VPWR VPWR U$$4010/A
+ sky130_fd_sc_hd__a22o_1
Xfanout574 U$$2196/X VGND VGND VPWR VPWR U$$2282/A2 sky130_fd_sc_hd__buf_4
XFILLER_59_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout585 U$$2006/A2 VGND VGND VPWR VPWR U$$1964/A2 sky130_fd_sc_hd__buf_4
Xfanout596 U$$1891/A2 VGND VGND VPWR VPWR U$$1859/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3308 U$$3580/B1 U$$3390/A2 U$$4406/A1 U$$3390/B2 VGND VGND VPWR VPWR U$$3309/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3319 U$$3319/A U$$3341/B VGND VGND VPWR VPWR U$$3319/X sky130_fd_sc_hd__xor2_1
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2607 U$$2605/Y input32/X U$$2603/A U$$2606/X U$$2603/Y VGND VGND VPWR VPWR U$$2607/X
+ sky130_fd_sc_hd__a32o_4
XU$$2618 U$$2618/A U$$2662/B VGND VGND VPWR VPWR U$$2618/X sky130_fd_sc_hd__xor2_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2629 U$$2629/A1 U$$2667/A2 U$$2631/A1 U$$2667/B2 VGND VGND VPWR VPWR U$$2630/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1906 U$$1906/A U$$1910/B VGND VGND VPWR VPWR U$$1906/X sky130_fd_sc_hd__xor2_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1917 input20/X VGND VGND VPWR VPWR U$$1917/Y sky130_fd_sc_hd__inv_1
XU$$1928 U$$3022/B1 U$$1964/A2 U$$2887/B1 U$$1964/B2 VGND VGND VPWR VPWR U$$1929/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ _408_/CLK _403_/D VGND VGND VPWR VPWR _403_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1939 U$$1939/A U$$1971/B VGND VGND VPWR VPWR U$$1939/X sky130_fd_sc_hd__xor2_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ _353_/CLK _334_/D VGND VGND VPWR VPWR _334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_265_ _397_/CLK _265_/D VGND VGND VPWR VPWR _265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_196_ _328_/CLK _196_/D VGND VGND VPWR VPWR _196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_95_0 dadda_fa_3_95_0/A dadda_fa_3_95_0/B dadda_fa_3_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_0/B dadda_fa_4_95_1/CIN sky130_fd_sc_hd__fa_1
XU$$554_1909 VGND VGND VPWR VPWR U$$554_1909/HI U$$554/A1 sky130_fd_sc_hd__conb_1
XFILLER_115_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4510 U$$811/A1 U$$4388/X U$$4512/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4511/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_57_5 dadda_fa_2_57_5/A dadda_fa_2_57_5/B dadda_fa_2_57_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_2/A dadda_fa_4_57_0/A sky130_fd_sc_hd__fa_1
XFILLER_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$13 U$$13/A U$$9/B VGND VGND VPWR VPWR U$$13/X sky130_fd_sc_hd__xor2_1
XU$$24 U$$24/A1 U$$48/A2 U$$26/A1 U$$48/B2 VGND VGND VPWR VPWR U$$25/A sky130_fd_sc_hd__a22o_1
XFILLER_65_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$35 U$$35/A U$$77/B VGND VGND VPWR VPWR U$$35/X sky130_fd_sc_hd__xor2_1
XU$$3820 U$$3820/A U$$3828/B VGND VGND VPWR VPWR U$$3820/X sky130_fd_sc_hd__xor2_1
XU$$3831 U$$4240/B1 U$$3833/A2 U$$4107/A1 U$$3833/B2 VGND VGND VPWR VPWR U$$3832/A
+ sky130_fd_sc_hd__a22o_1
XU$$46 U$$46/A1 U$$8/A2 U$$48/A1 U$$8/B2 VGND VGND VPWR VPWR U$$47/A sky130_fd_sc_hd__a22o_1
XU$$57 U$$57/A U$$87/B VGND VGND VPWR VPWR U$$57/X sky130_fd_sc_hd__xor2_1
XFILLER_92_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3842 U$$3842/A1 U$$3924/A2 U$$3979/B1 U$$3924/B2 VGND VGND VPWR VPWR U$$3843/A
+ sky130_fd_sc_hd__a22o_1
XU$$3853 U$$3853/A U$$3867/B VGND VGND VPWR VPWR U$$3853/X sky130_fd_sc_hd__xor2_1
XU$$3864 U$$3999/B1 U$$3892/A2 U$$4001/B1 U$$3892/B2 VGND VGND VPWR VPWR U$$3865/A
+ sky130_fd_sc_hd__a22o_1
XU$$68 U$$68/A1 U$$86/A2 U$$70/A1 U$$86/B2 VGND VGND VPWR VPWR U$$69/A sky130_fd_sc_hd__a22o_1
XU$$79 U$$79/A U$$81/B VGND VGND VPWR VPWR U$$79/X sky130_fd_sc_hd__xor2_1
XU$$3875 U$$3875/A U$$3925/B VGND VGND VPWR VPWR U$$3875/X sky130_fd_sc_hd__xor2_1
XU$$3886 U$$4434/A1 U$$3906/A2 U$$4162/A1 U$$3906/B2 VGND VGND VPWR VPWR U$$3887/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3897 U$$3897/A U$$3907/B VGND VGND VPWR VPWR U$$3897/X sky130_fd_sc_hd__xor2_1
XFILLER_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_96_0_1943 VGND VGND VPWR VPWR dadda_ha_1_96_0/A dadda_ha_1_96_0_1943/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_87_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_52_4 U$$1973/X U$$2106/X U$$2239/X VGND VGND VPWR VPWR dadda_fa_2_53_1/CIN
+ dadda_fa_2_52_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_45_3 U$$1294/X U$$1427/X U$$1560/X VGND VGND VPWR VPWR dadda_fa_2_46_3/A
+ dadda_fa_2_45_5/B sky130_fd_sc_hd__fa_1
XFILLER_55_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_22_2 dadda_fa_4_22_2/A dadda_fa_4_22_2/B dadda_fa_4_22_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_23_0/CIN dadda_fa_5_22_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_71_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_15_1 U$$702/X U$$835/X U$$968/X VGND VGND VPWR VPWR dadda_fa_5_16_0/B
+ dadda_fa_5_15_1/B sky130_fd_sc_hd__fa_1
XFILLER_52_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$1007 final_adder.U$$236/A final_adder.U$$737/X final_adder.U$$237/A2
+ VGND VGND VPWR VPWR final_adder.U$$1043/B sky130_fd_sc_hd__a21o_1
XFILLER_20_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1029 final_adder.U$$5/SUM final_adder.U$$1029/B VGND VGND VPWR VPWR
+ output340/A sky130_fd_sc_hd__xor2_1
XFILLER_165_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1303 fanout1309/X VGND VGND VPWR VPWR U$$3973/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1314 U$$3792/B VGND VGND VPWR VPWR U$$3790/B sky130_fd_sc_hd__buf_6
XFILLER_121_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1325 U$$955/B VGND VGND VPWR VPWR U$$907/B sky130_fd_sc_hd__buf_6
Xfanout1336 input49/X VGND VGND VPWR VPWR U$$3659/B sky130_fd_sc_hd__buf_4
XFILLER_66_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1347 input44/X VGND VGND VPWR VPWR U$$3341/B sky130_fd_sc_hd__buf_4
Xfanout1358 fanout1364/X VGND VGND VPWR VPWR U$$3288/A sky130_fd_sc_hd__buf_4
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1369 U$$3123/B VGND VGND VPWR VPWR U$$3077/B sky130_fd_sc_hd__buf_6
XFILLER_120_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout393 U$$952/A2 VGND VGND VPWR VPWR U$$902/A2 sky130_fd_sc_hd__clkbuf_8
XU$$3105 U$$3105/A U$$3107/B VGND VGND VPWR VPWR U$$3105/X sky130_fd_sc_hd__xor2_1
XFILLER_4_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3116 U$$4486/A1 U$$3118/A2 U$$4486/B1 U$$3118/B2 VGND VGND VPWR VPWR U$$3117/A
+ sky130_fd_sc_hd__a22o_1
XU$$3127 U$$3127/A U$$3150/A VGND VGND VPWR VPWR U$$3127/X sky130_fd_sc_hd__xor2_1
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3138 U$$3960/A1 U$$3144/A2 U$$3960/B1 U$$3144/B2 VGND VGND VPWR VPWR U$$3139/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2404 U$$2404/A U$$2408/B VGND VGND VPWR VPWR U$$2404/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3149 U$$3149/A U$$3150/A VGND VGND VPWR VPWR U$$3149/X sky130_fd_sc_hd__xor2_1
XU$$2415 U$$4196/A1 U$$2415/A2 U$$4196/B1 U$$2415/B2 VGND VGND VPWR VPWR U$$2416/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2426 U$$2426/A U$$2446/B VGND VGND VPWR VPWR U$$2426/X sky130_fd_sc_hd__xor2_1
XU$$2437 U$$2574/A1 U$$2443/A2 U$$2576/A1 U$$2443/B2 VGND VGND VPWR VPWR U$$2438/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2448 U$$2448/A U$$2456/B VGND VGND VPWR VPWR U$$2448/X sky130_fd_sc_hd__xor2_1
XU$$1703 U$$1703/A U$$1703/B VGND VGND VPWR VPWR U$$1703/X sky130_fd_sc_hd__xor2_1
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1714 U$$479/B1 U$$1720/A2 U$$346/A1 U$$1720/B2 VGND VGND VPWR VPWR U$$1715/A sky130_fd_sc_hd__a22o_1
XU$$2459 U$$952/A1 U$$2459/A2 U$$954/A1 U$$2459/B2 VGND VGND VPWR VPWR U$$2460/A sky130_fd_sc_hd__a22o_1
XU$$1725 U$$1725/A U$$1727/B VGND VGND VPWR VPWR U$$1725/X sky130_fd_sc_hd__xor2_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1736 U$$503/A1 U$$1774/A2 U$$505/A1 U$$1774/B2 VGND VGND VPWR VPWR U$$1737/A sky130_fd_sc_hd__a22o_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_973 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1747 U$$1747/A U$$1761/B VGND VGND VPWR VPWR U$$1747/X sky130_fd_sc_hd__xor2_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1758 U$$386/B1 U$$1758/A2 U$$253/A1 U$$1758/B2 VGND VGND VPWR VPWR U$$1759/A sky130_fd_sc_hd__a22o_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1769 U$$1769/A U$$1777/B VGND VGND VPWR VPWR U$$1769/X sky130_fd_sc_hd__xor2_1
XFILLER_42_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_317_ _321_/CLK _317_/D VGND VGND VPWR VPWR _317_/Q sky130_fd_sc_hd__dfxtp_1
Xinput13 a[20] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput24 a[30] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__dlymetal6s2s_1
X_248_ _377_/CLK _248_/D VGND VGND VPWR VPWR _248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput35 a[40] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
Xinput46 a[50] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__clkbuf_1
Xinput57 a[60] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_1
Xinput68 b[12] VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__clkbuf_4
X_179_ _328_/CLK _179_/D VGND VGND VPWR VPWR _179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput79 b[22] VGND VGND VPWR VPWR input79/X sky130_fd_sc_hd__buf_4
XFILLER_143_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_62_3 dadda_fa_2_62_3/A dadda_fa_2_62_3/B dadda_fa_2_62_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_1/B dadda_fa_3_62_3/B sky130_fd_sc_hd__fa_1
XFILLER_97_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_55_2 dadda_fa_2_55_2/A dadda_fa_2_55_2/B dadda_fa_2_55_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_1/A dadda_fa_3_55_3/A sky130_fd_sc_hd__fa_1
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_32_1 dadda_fa_5_32_1/A dadda_fa_5_32_1/B dadda_fa_5_32_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_33_0/B dadda_fa_7_32_0/A sky130_fd_sc_hd__fa_1
XU$$4340 U$$4340/A U$$4360/B VGND VGND VPWR VPWR U$$4340/X sky130_fd_sc_hd__xor2_1
XU$$4351 U$$4486/B1 U$$4373/A2 U$$4353/A1 U$$4373/B2 VGND VGND VPWR VPWR U$$4352/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_48_1 input199/X dadda_fa_2_48_1/B dadda_fa_2_48_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_49_0/CIN dadda_fa_3_48_2/CIN sky130_fd_sc_hd__fa_1
XU$$4362 U$$4362/A U$$4368/B VGND VGND VPWR VPWR U$$4362/X sky130_fd_sc_hd__xor2_1
XFILLER_53_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4373 U$$4508/B1 U$$4373/A2 U$$4375/A1 U$$4373/B2 VGND VGND VPWR VPWR U$$4374/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4384 U$$4384/A VGND VGND VPWR VPWR U$$4384/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_5_25_0 dadda_fa_5_25_0/A dadda_fa_5_25_0/B dadda_fa_5_25_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_26_0/A dadda_fa_6_25_0/CIN sky130_fd_sc_hd__fa_1
XU$$4395 U$$4395/A U$$4395/B VGND VGND VPWR VPWR U$$4395/X sky130_fd_sc_hd__xor2_1
XU$$3650 U$$3650/A1 U$$3696/A2 U$$3650/B1 U$$3696/B2 VGND VGND VPWR VPWR U$$3651/A
+ sky130_fd_sc_hd__a22o_1
XU$$3661 U$$3661/A U$$3681/B VGND VGND VPWR VPWR U$$3661/X sky130_fd_sc_hd__xor2_1
XFILLER_92_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3672 U$$4492/B1 U$$3682/A2 U$$4359/A1 U$$3682/B2 VGND VGND VPWR VPWR U$$3673/A
+ sky130_fd_sc_hd__a22o_1
XU$$3683 U$$3683/A U$$3695/B VGND VGND VPWR VPWR U$$3683/X sky130_fd_sc_hd__xor2_1
XU$$3694 U$$4240/B1 U$$3696/A2 U$$4107/A1 U$$3696/B2 VGND VGND VPWR VPWR U$$3695/A
+ sky130_fd_sc_hd__a22o_1
XU$$2960 U$$2960/A U$$2974/B VGND VGND VPWR VPWR U$$2960/X sky130_fd_sc_hd__xor2_1
XU$$2971 U$$3106/B1 U$$2979/A2 U$$2973/A1 U$$2979/B2 VGND VGND VPWR VPWR U$$2972/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2982 U$$2982/A U$$2986/B VGND VGND VPWR VPWR U$$2982/X sky130_fd_sc_hd__xor2_1
XU$$2993 U$$251/B1 U$$3005/A2 U$$2993/B1 U$$3005/B2 VGND VGND VPWR VPWR U$$2994/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4397_1846 VGND VGND VPWR VPWR U$$4397_1846/HI U$$4397/B sky130_fd_sc_hd__conb_1
XFILLER_20_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_37_1 U$$480/X U$$613/X VGND VGND VPWR VPWR dadda_fa_2_38_5/A dadda_fa_3_37_0/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$911 final_adder.U$$140/A final_adder.U$$849/X final_adder.U$$911/B1
+ VGND VGND VPWR VPWR final_adder.U$$911/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$933 final_adder.U$$162/A final_adder.U$$871/X final_adder.U$$933/B1
+ VGND VGND VPWR VPWR final_adder.U$$933/X sky130_fd_sc_hd__a21o_1
XFILLER_169_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_50_1 U$$506/X U$$639/X U$$772/X VGND VGND VPWR VPWR dadda_fa_2_51_0/CIN
+ dadda_fa_2_50_3/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$955 final_adder.U$$184/A final_adder.U$$893/X final_adder.U$$955/B1
+ VGND VGND VPWR VPWR final_adder.U$$955/X sky130_fd_sc_hd__a21o_1
XU$$805 U$$805/A1 U$$807/A2 U$$805/B1 U$$807/B2 VGND VGND VPWR VPWR U$$806/A sky130_fd_sc_hd__a22o_1
XFILLER_113_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$977 final_adder.U$$206/A final_adder.U$$819/X final_adder.U$$977/B1
+ VGND VGND VPWR VPWR final_adder.U$$977/X sky130_fd_sc_hd__a21o_1
Xclkbuf_2_2__f_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _388_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$816 U$$816/A U$$820/B VGND VGND VPWR VPWR U$$816/X sky130_fd_sc_hd__xor2_1
XU$$827 U$$825/B U$$822/A input4/X U$$822/Y VGND VGND VPWR VPWR U$$827/X sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_43_0 U$$93/X U$$226/X U$$359/X VGND VGND VPWR VPWR dadda_fa_2_44_2/CIN
+ dadda_fa_2_43_4/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$999 final_adder.U$$228/A final_adder.U$$729/X final_adder.U$$999/B1
+ VGND VGND VPWR VPWR final_adder.U$$999/X sky130_fd_sc_hd__a21o_1
XFILLER_83_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$838 U$$973/B1 U$$904/A2 U$$840/A1 U$$904/B2 VGND VGND VPWR VPWR U$$839/A sky130_fd_sc_hd__a22o_1
XU$$849 U$$849/A U$$907/B VGND VGND VPWR VPWR U$$849/X sky130_fd_sc_hd__xor2_1
XFILLER_43_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_72_2 dadda_fa_3_72_2/A dadda_fa_3_72_2/B dadda_fa_3_72_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_1/A dadda_fa_4_72_2/B sky130_fd_sc_hd__fa_1
XFILLER_105_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1100 U$$3618/A1 VGND VGND VPWR VPWR U$$4440/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_152_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_65_1 dadda_fa_3_65_1/A dadda_fa_3_65_1/B dadda_fa_3_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_0/CIN dadda_fa_4_65_2/A sky130_fd_sc_hd__fa_1
Xfanout1111 U$$735/B1 VGND VGND VPWR VPWR U$$52/A1 sky130_fd_sc_hd__buf_4
Xfanout1122 U$$3610/B1 VGND VGND VPWR VPWR U$$872/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_152_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1133 input77/X VGND VGND VPWR VPWR U$$3884/A1 sky130_fd_sc_hd__buf_4
XFILLER_152_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1144 input75/X VGND VGND VPWR VPWR U$$2923/A1 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_6_42_0 dadda_fa_6_42_0/A dadda_fa_6_42_0/B dadda_fa_6_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_43_0/B dadda_fa_7_42_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_58_0 dadda_fa_3_58_0/A dadda_fa_3_58_0/B dadda_fa_3_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_0/B dadda_fa_4_58_1/CIN sky130_fd_sc_hd__fa_1
Xfanout1155 U$$316/B1 VGND VGND VPWR VPWR U$$44/A1 sky130_fd_sc_hd__buf_4
XFILLER_121_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1166 U$$4424/B1 VGND VGND VPWR VPWR U$$4152/A1 sky130_fd_sc_hd__buf_6
Xfanout1177 U$$3189/A1 VGND VGND VPWR VPWR U$$997/A1 sky130_fd_sc_hd__buf_4
Xfanout1188 input70/X VGND VGND VPWR VPWR U$$3870/B1 sky130_fd_sc_hd__buf_6
Xfanout1199 U$$1088/B VGND VGND VPWR VPWR U$$982/B sky130_fd_sc_hd__buf_6
XFILLER_93_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2201 U$$2201/A U$$2253/B VGND VGND VPWR VPWR U$$2201/X sky130_fd_sc_hd__xor2_1
XFILLER_90_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2212 U$$4404/A1 U$$2252/A2 U$$2897/B1 U$$2252/B2 VGND VGND VPWR VPWR U$$2213/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_101_2 dadda_fa_4_101_2/A dadda_fa_4_101_2/B dadda_fa_4_101_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_102_0/CIN dadda_fa_5_101_1/CIN sky130_fd_sc_hd__fa_1
XU$$2223 U$$2223/A U$$2231/B VGND VGND VPWR VPWR U$$2223/X sky130_fd_sc_hd__xor2_1
XFILLER_90_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2234 U$$40/B1 U$$2252/A2 U$$316/B1 U$$2252/B2 VGND VGND VPWR VPWR U$$2235/A sky130_fd_sc_hd__a22o_1
XU$$1500 U$$539/B1 U$$1502/A2 U$$406/A1 U$$1502/B2 VGND VGND VPWR VPWR U$$1501/A sky130_fd_sc_hd__a22o_1
XFILLER_62_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2245 U$$2245/A U$$2283/B VGND VGND VPWR VPWR U$$2245/X sky130_fd_sc_hd__xor2_1
XU$$1511 U$$1509/Y input15/X U$$1507/A U$$1510/X U$$1507/Y VGND VGND VPWR VPWR U$$1511/X
+ sky130_fd_sc_hd__a32o_1
XU$$2256 U$$2665/B1 U$$2272/A2 U$$66/A1 U$$2272/B2 VGND VGND VPWR VPWR U$$2257/A sky130_fd_sc_hd__a22o_1
XU$$1522 U$$1522/A U$$1564/B VGND VGND VPWR VPWR U$$1522/X sky130_fd_sc_hd__xor2_1
XU$$2267 U$$2267/A U$$2301/B VGND VGND VPWR VPWR U$$2267/X sky130_fd_sc_hd__xor2_1
XU$$1533 U$$2629/A1 U$$1575/A2 U$$2631/A1 U$$1575/B2 VGND VGND VPWR VPWR U$$1534/A
+ sky130_fd_sc_hd__a22o_1
XU$$2278 U$$906/B1 U$$2282/A2 U$$773/A1 U$$2282/B2 VGND VGND VPWR VPWR U$$2279/A sky130_fd_sc_hd__a22o_1
XFILLER_62_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1544 U$$1544/A U$$1584/B VGND VGND VPWR VPWR U$$1544/X sky130_fd_sc_hd__xor2_1
XU$$2289 U$$2289/A U$$2327/B VGND VGND VPWR VPWR U$$2289/X sky130_fd_sc_hd__xor2_1
XFILLER_31_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1555 U$$596/A1 U$$1563/A2 U$$596/B1 U$$1563/B2 VGND VGND VPWR VPWR U$$1556/A sky130_fd_sc_hd__a22o_1
XU$$1566 U$$1566/A U$$1568/B VGND VGND VPWR VPWR U$$1566/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_116_0 dadda_ha_3_116_0/A U$$3697/X VGND VGND VPWR VPWR dadda_fa_4_117_2/CIN
+ dadda_ha_3_116_0/SUM sky130_fd_sc_hd__ha_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1577 U$$481/A1 U$$1587/A2 U$$72/A1 U$$1587/B2 VGND VGND VPWR VPWR U$$1578/A sky130_fd_sc_hd__a22o_1
XFILLER_15_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1588 U$$1588/A U$$1618/B VGND VGND VPWR VPWR U$$1588/X sky130_fd_sc_hd__xor2_1
XU$$1599 U$$3106/A1 U$$1635/A2 U$$3106/B1 U$$1635/B2 VGND VGND VPWR VPWR U$$1600/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_115_0 dadda_fa_7_115_0/A dadda_fa_7_115_0/B dadda_fa_7_115_0/CIN VGND
+ VGND VPWR VPWR _412_/D _283_/D sky130_fd_sc_hd__fa_1
XFILLER_147_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_0 dadda_fa_2_60_0/A dadda_fa_2_60_0/B dadda_fa_2_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_0/B dadda_fa_3_60_2/B sky130_fd_sc_hd__fa_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$207 final_adder.U$$206/B final_adder.U$$977/B1 final_adder.U$$207/B1
+ VGND VGND VPWR VPWR final_adder.U$$207/X sky130_fd_sc_hd__a21o_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$218 final_adder.U$$218/A final_adder.U$$218/B VGND VGND VPWR VPWR
+ final_adder.U$$346/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$229 final_adder.U$$228/B final_adder.U$$999/B1 final_adder.U$$229/B1
+ VGND VGND VPWR VPWR final_adder.U$$229/X sky130_fd_sc_hd__a21o_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4170 U$$4307/A1 U$$4174/A2 U$$4307/B1 U$$4174/B2 VGND VGND VPWR VPWR U$$4171/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4181 U$$4181/A U$$4231/B VGND VGND VPWR VPWR U$$4181/X sky130_fd_sc_hd__xor2_1
XU$$4192 U$$4464/B1 U$$4224/A2 U$$4331/A1 U$$4224/B2 VGND VGND VPWR VPWR U$$4193/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3480 U$$3480/A U$$3524/B VGND VGND VPWR VPWR U$$3480/X sky130_fd_sc_hd__xor2_1
XU$$3491 U$$3628/A1 U$$3505/A2 U$$3628/B1 U$$3505/B2 VGND VGND VPWR VPWR U$$3492/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2790 U$$3338/A1 U$$2798/A2 U$$735/B1 U$$2798/B2 VGND VGND VPWR VPWR U$$2791/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_82_1 dadda_fa_4_82_1/A dadda_fa_4_82_1/B dadda_fa_4_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_83_0/B dadda_fa_5_82_1/B sky130_fd_sc_hd__fa_1
XFILLER_134_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_75_0 dadda_fa_4_75_0/A dadda_fa_4_75_0/B dadda_fa_4_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_76_0/A dadda_fa_5_75_1/A sky130_fd_sc_hd__fa_1
XFILLER_0_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput203 c[51] VGND VGND VPWR VPWR input203/X sky130_fd_sc_hd__buf_2
XFILLER_88_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4451_1873 VGND VGND VPWR VPWR U$$4451_1873/HI U$$4451/B sky130_fd_sc_hd__conb_1
Xinput214 c[61] VGND VGND VPWR VPWR input214/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput225 c[71] VGND VGND VPWR VPWR input225/X sky130_fd_sc_hd__clkbuf_2
Xinput236 c[81] VGND VGND VPWR VPWR input236/X sky130_fd_sc_hd__clkbuf_2
Xinput247 c[91] VGND VGND VPWR VPWR input247/X sky130_fd_sc_hd__buf_2
XFILLER_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$741 final_adder.U$$740/B final_adder.U$$661/X final_adder.U$$629/X
+ VGND VGND VPWR VPWR final_adder.U$$741/X sky130_fd_sc_hd__a21o_1
XFILLER_84_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$752 final_adder.U$$784/B final_adder.U$$752/B VGND VGND VPWR VPWR
+ final_adder.U$$752/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$763 final_adder.U$$762/B final_adder.U$$683/X final_adder.U$$651/X
+ VGND VGND VPWR VPWR final_adder.U$$763/X sky130_fd_sc_hd__a21o_1
XFILLER_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$602 U$$602/A1 U$$636/A2 U$$56/A1 U$$636/B2 VGND VGND VPWR VPWR U$$603/A sky130_fd_sc_hd__a22o_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$774 final_adder.U$$774/A final_adder.U$$774/B VGND VGND VPWR VPWR
+ final_adder.U$$774/X sky130_fd_sc_hd__and2_1
XFILLER_44_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$613 U$$613/A U$$643/B VGND VGND VPWR VPWR U$$613/X sky130_fd_sc_hd__xor2_1
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$785 final_adder.U$$784/B final_adder.U$$705/X final_adder.U$$673/X
+ VGND VGND VPWR VPWR final_adder.U$$785/X sky130_fd_sc_hd__a21o_1
XU$$624 U$$898/A1 U$$630/A2 U$$900/A1 U$$630/B2 VGND VGND VPWR VPWR U$$625/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$796 final_adder.U$$796/A final_adder.U$$796/B VGND VGND VPWR VPWR
+ final_adder.U$$796/X sky130_fd_sc_hd__and2_1
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$635 U$$635/A U$$637/B VGND VGND VPWR VPWR U$$635/X sky130_fd_sc_hd__xor2_1
XU$$646 U$$783/A1 U$$682/A2 U$$783/B1 U$$682/B2 VGND VGND VPWR VPWR U$$647/A sky130_fd_sc_hd__a22o_1
XU$$657 U$$657/A U$$669/B VGND VGND VPWR VPWR U$$657/X sky130_fd_sc_hd__xor2_1
XFILLER_83_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$668 U$$805/A1 U$$674/A2 U$$805/B1 U$$674/B2 VGND VGND VPWR VPWR U$$669/A sky130_fd_sc_hd__a22o_1
XFILLER_140_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$679 U$$679/A U$$684/A VGND VGND VPWR VPWR U$$679/X sky130_fd_sc_hd__xor2_1
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_889 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_32_4 U$$1667/X U$$1800/X U$$1933/X VGND VGND VPWR VPWR dadda_fa_3_33_1/CIN
+ dadda_fa_3_32_3/CIN sky130_fd_sc_hd__fa_1
XU$$2020 U$$4486/A1 U$$2052/A2 U$$4486/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2021/A
+ sky130_fd_sc_hd__a22o_1
XU$$2031 U$$2031/A U$$2031/B VGND VGND VPWR VPWR U$$2031/X sky130_fd_sc_hd__xor2_1
XFILLER_74_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2042 U$$2042/A1 U$$2044/A2 U$$2179/B1 U$$2044/B2 VGND VGND VPWR VPWR U$$2043/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2053 U$$2053/A U$$2053/B VGND VGND VPWR VPWR U$$2053/X sky130_fd_sc_hd__xor2_1
XFILLER_35_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2064 U$$2064/A U$$2096/B VGND VGND VPWR VPWR U$$2064/X sky130_fd_sc_hd__xor2_1
XU$$1330 U$$1330/A U$$1364/B VGND VGND VPWR VPWR U$$1330/X sky130_fd_sc_hd__xor2_1
XU$$2075 U$$840/B1 U$$2107/A2 U$$707/A1 U$$2107/B2 VGND VGND VPWR VPWR U$$2076/A sky130_fd_sc_hd__a22o_1
XU$$2086 U$$2086/A U$$2096/B VGND VGND VPWR VPWR U$$2086/X sky130_fd_sc_hd__xor2_1
XU$$1341 U$$930/A1 U$$1361/A2 U$$2711/B1 U$$1361/B2 VGND VGND VPWR VPWR U$$1342/A
+ sky130_fd_sc_hd__a22o_1
XU$$2097 U$$999/B1 U$$2097/A2 U$$866/A1 U$$2097/B2 VGND VGND VPWR VPWR U$$2098/A sky130_fd_sc_hd__a22o_1
XU$$1352 U$$1352/A U$$1358/B VGND VGND VPWR VPWR U$$1352/X sky130_fd_sc_hd__xor2_1
XU$$1363 U$$539/B1 U$$1367/A2 U$$406/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1364/A sky130_fd_sc_hd__a22o_1
XFILLER_149_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1374 U$$1372/Y input13/X U$$1370/A U$$1373/X U$$1370/Y VGND VGND VPWR VPWR U$$1374/X
+ sky130_fd_sc_hd__a32o_1
XU$$1385 U$$1385/A U$$1427/B VGND VGND VPWR VPWR U$$1385/X sky130_fd_sc_hd__xor2_1
XU$$1396 U$$983/B1 U$$1432/A2 U$$850/A1 U$$1432/B2 VGND VGND VPWR VPWR U$$1397/A sky130_fd_sc_hd__a22o_1
XFILLER_117_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_92_0 dadda_fa_5_92_0/A dadda_fa_5_92_0/B dadda_fa_5_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_93_0/A dadda_fa_6_92_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_128_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout904 U$$1194/B2 VGND VGND VPWR VPWR U$$1164/B2 sky130_fd_sc_hd__buf_4
XFILLER_143_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout915 U$$48/B2 VGND VGND VPWR VPWR U$$8/B2 sky130_fd_sc_hd__buf_2
Xdadda_fa_1_77_6 U$$3752/X U$$3885/X U$$4018/X VGND VGND VPWR VPWR dadda_fa_2_78_2/B
+ dadda_fa_2_77_5/B sky130_fd_sc_hd__fa_1
Xfanout926 U$$4502/B2 VGND VGND VPWR VPWR U$$4488/B2 sky130_fd_sc_hd__clkbuf_4
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout937 fanout938/X VGND VGND VPWR VPWR U$$910/A1 sky130_fd_sc_hd__buf_4
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout948 input98/X VGND VGND VPWR VPWR U$$4398/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_97_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout959 fanout966/X VGND VGND VPWR VPWR U$$84/A1 sky130_fd_sc_hd__buf_2
XFILLER_38_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$70 _366_/Q _238_/Q VGND VGND VPWR VPWR final_adder.U$$955/B1 final_adder.U$$184/A
+ sky130_fd_sc_hd__ha_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$81 _377_/Q _249_/Q VGND VGND VPWR VPWR final_adder.U$$175/B1 final_adder.U$$174/B
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$92 _388_/Q _260_/Q VGND VGND VPWR VPWR final_adder.U$$933/B1 final_adder.U$$162/A
+ sky130_fd_sc_hd__ha_1
XU$$4481_1888 VGND VGND VPWR VPWR U$$4481_1888/HI U$$4481/B sky130_fd_sc_hd__conb_1
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_101_1 input131/X dadda_fa_3_101_1/B dadda_fa_3_101_1/CIN VGND VGND VPWR
+ VPWR dadda_fa_4_102_0/CIN dadda_fa_4_101_2/A sky130_fd_sc_hd__fa_1
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_122_0 dadda_fa_6_122_0/A dadda_fa_6_122_0/B dadda_fa_6_122_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_123_0/B dadda_fa_7_122_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_65_4 U$$1733/X U$$1866/X U$$1999/X VGND VGND VPWR VPWR dadda_fa_1_66_6/CIN
+ dadda_fa_1_65_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_42_3 dadda_fa_3_42_3/A dadda_fa_3_42_3/B dadda_fa_3_42_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_1/B dadda_fa_4_42_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$560 final_adder.U$$568/B final_adder.U$$560/B VGND VGND VPWR VPWR
+ final_adder.U$$680/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$571 final_adder.U$$570/B final_adder.U$$455/X final_adder.U$$447/X
+ VGND VGND VPWR VPWR final_adder.U$$571/X sky130_fd_sc_hd__a21o_1
XFILLER_29_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$410 U$$410/A VGND VGND VPWR VPWR U$$410/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$582 final_adder.U$$590/B final_adder.U$$582/B VGND VGND VPWR VPWR
+ final_adder.U$$702/B sky130_fd_sc_hd__and2_1
XFILLER_57_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_35_2 dadda_fa_3_35_2/A dadda_fa_3_35_2/B dadda_fa_3_35_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_1/A dadda_fa_4_35_2/B sky130_fd_sc_hd__fa_1
XU$$421 U$$10/A1 U$$447/A2 U$$12/A1 U$$447/B2 VGND VGND VPWR VPWR U$$422/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$593 final_adder.U$$592/B final_adder.U$$477/X final_adder.U$$469/X
+ VGND VGND VPWR VPWR final_adder.U$$593/X sky130_fd_sc_hd__a21o_1
XU$$432 U$$432/A U$$448/B VGND VGND VPWR VPWR U$$432/X sky130_fd_sc_hd__xor2_1
XFILLER_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$443 U$$443/A1 U$$505/A2 U$$34/A1 U$$505/B2 VGND VGND VPWR VPWR U$$444/A sky130_fd_sc_hd__a22o_1
XFILLER_44_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$454 U$$454/A U$$504/B VGND VGND VPWR VPWR U$$454/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_28_1 U$$1925/X U$$1963/B input177/X VGND VGND VPWR VPWR dadda_fa_4_29_0/CIN
+ dadda_fa_4_28_2/A sky130_fd_sc_hd__fa_1
XU$$465 U$$465/A1 U$$501/A2 U$$465/B1 U$$501/B2 VGND VGND VPWR VPWR U$$466/A sky130_fd_sc_hd__a22o_1
XFILLER_60_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$476 U$$476/A U$$480/B VGND VGND VPWR VPWR U$$476/X sky130_fd_sc_hd__xor2_1
XU$$487 U$$487/A1 U$$501/A2 U$$487/B1 U$$501/B2 VGND VGND VPWR VPWR U$$488/A sky130_fd_sc_hd__a22o_1
XU$$498 U$$498/A U$$498/B VGND VGND VPWR VPWR U$$498/X sky130_fd_sc_hd__xor2_1
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_87_5 dadda_fa_2_87_5/A dadda_fa_2_87_5/B dadda_fa_2_87_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_88_2/A dadda_fa_4_87_0/A sky130_fd_sc_hd__fa_2
XFILLER_119_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_30_1 U$$466/X U$$599/X U$$732/X VGND VGND VPWR VPWR dadda_fa_3_31_1/B
+ dadda_fa_3_30_3/A sky130_fd_sc_hd__fa_1
XFILLER_63_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1160 U$$64/A1 U$$1164/A2 U$$64/B1 U$$1164/B2 VGND VGND VPWR VPWR U$$1161/A sky130_fd_sc_hd__a22o_1
XU$$1171 U$$1171/A U$$1171/B VGND VGND VPWR VPWR U$$1171/X sky130_fd_sc_hd__xor2_1
XU$$1182 U$$906/B1 U$$1218/A2 U$$773/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1183/A sky130_fd_sc_hd__a22o_1
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1193 U$$1193/A U$$1195/B VGND VGND VPWR VPWR U$$1193/X sky130_fd_sc_hd__xor2_1
XFILLER_149_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_117_1 dadda_fa_5_117_1/A dadda_fa_5_117_1/B dadda_fa_5_117_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_118_0/B dadda_fa_7_117_0/A sky130_fd_sc_hd__fa_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_82_4 U$$2831/X U$$2964/X U$$3097/X VGND VGND VPWR VPWR dadda_fa_2_83_2/CIN
+ dadda_fa_2_82_5/A sky130_fd_sc_hd__fa_1
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout701 U$$4244/B2 VGND VGND VPWR VPWR U$$4158/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout712 U$$3978/X VGND VGND VPWR VPWR U$$4043/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout723 U$$3966/B2 VGND VGND VPWR VPWR U$$3948/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_75_3 U$$2817/X U$$2950/X U$$3083/X VGND VGND VPWR VPWR dadda_fa_2_76_1/B
+ dadda_fa_2_75_4/B sky130_fd_sc_hd__fa_1
Xfanout734 U$$3704/X VGND VGND VPWR VPWR U$$3833/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout745 U$$3473/B2 VGND VGND VPWR VPWR U$$3511/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_52_2 dadda_fa_4_52_2/A dadda_fa_4_52_2/B dadda_fa_4_52_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_53_0/CIN dadda_fa_5_52_1/CIN sky130_fd_sc_hd__fa_1
Xfanout756 U$$3306/B2 VGND VGND VPWR VPWR U$$3390/B2 sky130_fd_sc_hd__buf_6
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_2 U$$3335/X U$$3468/X U$$3601/X VGND VGND VPWR VPWR dadda_fa_2_69_1/A
+ dadda_fa_2_68_4/A sky130_fd_sc_hd__fa_1
Xfanout767 U$$3251/B2 VGND VGND VPWR VPWR U$$3285/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout778 U$$3019/X VGND VGND VPWR VPWR U$$3118/B2 sky130_fd_sc_hd__buf_4
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout789 U$$408/B2 VGND VGND VPWR VPWR U$$406/B2 sky130_fd_sc_hd__buf_4
XFILLER_74_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_45_1 dadda_fa_4_45_1/A dadda_fa_4_45_1/B dadda_fa_4_45_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_46_0/B dadda_fa_5_45_1/B sky130_fd_sc_hd__fa_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_22_0 dadda_fa_7_22_0/A dadda_fa_7_22_0/B dadda_fa_7_22_0/CIN VGND VGND
+ VPWR VPWR _319_/D _190_/D sky130_fd_sc_hd__fa_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_38_0 dadda_fa_4_38_0/A dadda_fa_4_38_0/B dadda_fa_4_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_39_0/A dadda_fa_5_38_1/A sky130_fd_sc_hd__fa_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ _353_/CLK _350_/D VGND VGND VPWR VPWR _350_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_281_ _416_/CLK _281_/D VGND VGND VPWR VPWR _281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_0_57_2 U$$919/X U$$1052/X VGND VGND VPWR VPWR dadda_fa_1_58_7/CIN dadda_fa_2_57_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_70_2 U$$1211/X U$$1344/X U$$1477/X VGND VGND VPWR VPWR dadda_fa_1_71_7/A
+ dadda_fa_1_70_8/B sky130_fd_sc_hd__fa_1
XFILLER_65_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_63_1 U$$532/X U$$665/X U$$798/X VGND VGND VPWR VPWR dadda_fa_1_64_5/CIN
+ dadda_fa_1_63_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_40_0 dadda_fa_3_40_0/A dadda_fa_3_40_0/B dadda_fa_3_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_0/B dadda_fa_4_40_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_56_0 U$$119/X U$$252/X U$$385/X VGND VGND VPWR VPWR dadda_fa_1_57_7/B
+ dadda_fa_1_56_8/B sky130_fd_sc_hd__fa_1
XFILLER_64_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$390 final_adder.U$$394/B final_adder.U$$390/B VGND VGND VPWR VPWR
+ final_adder.U$$514/B sky130_fd_sc_hd__and2_1
XFILLER_18_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$240 U$$240/A U$$254/B VGND VGND VPWR VPWR U$$240/X sky130_fd_sc_hd__xor2_1
XU$$251 U$$251/A1 U$$253/A2 U$$251/B1 U$$253/B2 VGND VGND VPWR VPWR U$$252/A sky130_fd_sc_hd__a22o_1
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$262 U$$262/A U$$273/A VGND VGND VPWR VPWR U$$262/X sky130_fd_sc_hd__xor2_1
XU$$273 U$$273/A VGND VGND VPWR VPWR U$$273/Y sky130_fd_sc_hd__inv_1
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$284 U$$10/A1 U$$312/A2 U$$12/A1 U$$312/B2 VGND VGND VPWR VPWR U$$285/A sky130_fd_sc_hd__a22o_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$295 U$$295/A U$$347/B VGND VGND VPWR VPWR U$$295/X sky130_fd_sc_hd__xor2_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1 U$$1/A VGND VGND VPWR VPWR U$$3/B sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$9 _305_/Q _177_/Q VGND VGND VPWR VPWR final_adder.U$$9/COUT final_adder.U$$9/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput304 output304/A VGND VGND VPWR VPWR o[27] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_3 U$$4181/X U$$4314/X U$$4447/X VGND VGND VPWR VPWR dadda_fa_3_93_1/B
+ dadda_fa_3_92_3/B sky130_fd_sc_hd__fa_1
Xoutput315 output315/A VGND VGND VPWR VPWR o[37] sky130_fd_sc_hd__buf_2
Xoutput326 output326/A VGND VGND VPWR VPWR o[47] sky130_fd_sc_hd__buf_2
Xoutput337 output337/A VGND VGND VPWR VPWR o[57] sky130_fd_sc_hd__buf_2
XFILLER_114_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_85_2 dadda_fa_2_85_2/A dadda_fa_2_85_2/B dadda_fa_2_85_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_1/A dadda_fa_3_85_3/A sky130_fd_sc_hd__fa_1
Xoutput348 output348/A VGND VGND VPWR VPWR o[67] sky130_fd_sc_hd__buf_2
Xoutput359 output359/A VGND VGND VPWR VPWR o[77] sky130_fd_sc_hd__buf_2
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_62_1 dadda_fa_5_62_1/A dadda_fa_5_62_1/B dadda_fa_5_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_63_0/B dadda_fa_7_62_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_78_1 dadda_fa_2_78_1/A dadda_fa_2_78_1/B dadda_fa_2_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_0/CIN dadda_fa_3_78_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_55_0 dadda_fa_5_55_0/A dadda_fa_5_55_0/B dadda_fa_5_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_56_0/A dadda_fa_6_55_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_54_8 input206/X dadda_fa_1_54_8/B dadda_fa_1_54_8/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_55_3/A dadda_fa_3_54_0/A sky130_fd_sc_hd__fa_1
XFILLER_95_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_101_0 U$$2602/Y U$$2736/X U$$2869/X VGND VGND VPWR VPWR dadda_fa_3_102_1/CIN
+ dadda_fa_3_101_3/A sky130_fd_sc_hd__fa_1
XFILLER_36_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_80_1 U$$1497/X U$$1630/X U$$1763/X VGND VGND VPWR VPWR dadda_fa_2_81_1/A
+ dadda_fa_2_80_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1507 U$$985/A1 VGND VGND VPWR VPWR U$$2629/A1 sky130_fd_sc_hd__buf_4
Xfanout520 U$$2937/A2 VGND VGND VPWR VPWR U$$2929/A2 sky130_fd_sc_hd__buf_4
Xfanout1518 input127/X VGND VGND VPWR VPWR U$$4271/A1 sky130_fd_sc_hd__buf_4
XFILLER_104_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_73_0 U$$1882/X U$$2015/X U$$2148/X VGND VGND VPWR VPWR dadda_fa_2_74_0/B
+ dadda_fa_2_73_3/B sky130_fd_sc_hd__fa_1
Xfanout531 U$$278/X VGND VGND VPWR VPWR U$$408/A2 sky130_fd_sc_hd__buf_4
Xfanout1529 U$$4406/A1 VGND VGND VPWR VPWR U$$707/A1 sky130_fd_sc_hd__buf_4
Xfanout542 U$$2874/A2 VGND VGND VPWR VPWR U$$2872/A2 sky130_fd_sc_hd__buf_4
XFILLER_76_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout553 U$$2540/A2 VGND VGND VPWR VPWR U$$2532/A2 sky130_fd_sc_hd__buf_4
Xfanout564 U$$2445/A2 VGND VGND VPWR VPWR U$$2443/A2 sky130_fd_sc_hd__buf_6
Xfanout575 U$$2320/A2 VGND VGND VPWR VPWR U$$2310/A2 sky130_fd_sc_hd__buf_6
Xfanout586 U$$2022/A2 VGND VGND VPWR VPWR U$$2006/A2 sky130_fd_sc_hd__buf_4
XFILLER_74_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout597 U$$1881/A2 VGND VGND VPWR VPWR U$$1841/A2 sky130_fd_sc_hd__buf_6
XFILLER_74_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3309 U$$3309/A U$$3349/B VGND VGND VPWR VPWR U$$3309/X sky130_fd_sc_hd__xor2_1
XFILLER_58_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2608 U$$2606/B U$$2603/A input32/X U$$2603/Y VGND VGND VPWR VPWR U$$2608/X sky130_fd_sc_hd__a22o_4
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2619 U$$2891/B1 U$$2665/A2 U$$2758/A1 U$$2665/B2 VGND VGND VPWR VPWR U$$2620/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1907 U$$2179/B1 U$$1911/A2 U$$2183/A1 U$$1911/B2 VGND VGND VPWR VPWR U$$1908/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1918 U$$1918/A VGND VGND VPWR VPWR U$$1918/Y sky130_fd_sc_hd__inv_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_402_ _402_/CLK _402_/D VGND VGND VPWR VPWR _402_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1929 U$$1929/A U$$1963/B VGND VGND VPWR VPWR U$$1929/X sky130_fd_sc_hd__xor2_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_333_ _344_/CLK _333_/D VGND VGND VPWR VPWR _333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_264_ _397_/CLK _264_/D VGND VGND VPWR VPWR _264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_195_ _328_/CLK _195_/D VGND VGND VPWR VPWR _195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_95_1 dadda_fa_3_95_1/A dadda_fa_3_95_1/B dadda_fa_3_95_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_0/CIN dadda_fa_4_95_2/A sky130_fd_sc_hd__fa_1
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_72_0 dadda_fa_6_72_0/A dadda_fa_6_72_0/B dadda_fa_6_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_73_0/B dadda_fa_7_72_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_88_0 dadda_fa_3_88_0/A dadda_fa_3_88_0/B dadda_fa_3_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_0/B dadda_fa_4_88_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_2_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4500 U$$4500/A1 U$$4388/X U$$4502/A1 U$$4502/B2 VGND VGND VPWR VPWR U$$4501/A
+ sky130_fd_sc_hd__a22o_1
XU$$4511 U$$4511/A U$$4511/B VGND VGND VPWR VPWR U$$4511/X sky130_fd_sc_hd__xor2_1
XFILLER_49_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$14 U$$14/A1 U$$8/A2 U$$16/A1 U$$8/B2 VGND VGND VPWR VPWR U$$15/A sky130_fd_sc_hd__a22o_1
XU$$3810 U$$3810/A U$$3835/A VGND VGND VPWR VPWR U$$3810/X sky130_fd_sc_hd__xor2_1
XU$$25 U$$25/A U$$49/B VGND VGND VPWR VPWR U$$25/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_117_0 U$$3698/Y U$$3832/X U$$3965/X VGND VGND VPWR VPWR dadda_fa_5_118_0/A
+ dadda_fa_5_117_1/A sky130_fd_sc_hd__fa_1
XU$$3821 U$$4367/B1 U$$3829/A2 U$$4234/A1 U$$3829/B2 VGND VGND VPWR VPWR U$$3822/A
+ sky130_fd_sc_hd__a22o_1
XU$$36 U$$36/A1 U$$74/A2 U$$38/A1 U$$74/B2 VGND VGND VPWR VPWR U$$37/A sky130_fd_sc_hd__a22o_1
XU$$3832 U$$3832/A U$$3835/A VGND VGND VPWR VPWR U$$3832/X sky130_fd_sc_hd__xor2_1
XFILLER_65_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$47 U$$47/A U$$49/B VGND VGND VPWR VPWR U$$47/X sky130_fd_sc_hd__xor2_1
XU$$58 U$$58/A1 U$$96/A2 U$$60/A1 U$$96/B2 VGND VGND VPWR VPWR U$$59/A sky130_fd_sc_hd__a22o_1
XU$$3843 U$$3843/A U$$3925/B VGND VGND VPWR VPWR U$$3843/X sky130_fd_sc_hd__xor2_1
XU$$3854 U$$4400/B1 U$$3892/A2 U$$4265/B1 U$$3892/B2 VGND VGND VPWR VPWR U$$3855/A
+ sky130_fd_sc_hd__a22o_1
XU$$69 U$$69/A U$$87/B VGND VGND VPWR VPWR U$$69/X sky130_fd_sc_hd__xor2_1
XU$$3865 U$$3865/A U$$3867/B VGND VGND VPWR VPWR U$$3865/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_5_4_0 U$$15/X U$$148/X VGND VGND VPWR VPWR dadda_fa_6_5_0/CIN dadda_fa_7_4_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3876 U$$4150/A1 U$$3924/A2 U$$4152/A1 U$$3924/B2 VGND VGND VPWR VPWR U$$3877/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3887 U$$3887/A U$$3973/A VGND VGND VPWR VPWR U$$3887/X sky130_fd_sc_hd__xor2_1
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3898 U$$4307/B1 U$$3906/A2 U$$4174/A1 U$$3906/B2 VGND VGND VPWR VPWR U$$3899/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_90_0 U$$3246/X U$$3379/X U$$3512/X VGND VGND VPWR VPWR dadda_fa_3_91_0/B
+ dadda_fa_3_90_2/B sky130_fd_sc_hd__fa_1
XFILLER_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_46_6 U$$2493/X U$$2626/X VGND VGND VPWR VPWR dadda_fa_2_47_3/CIN dadda_fa_3_46_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_52_5 U$$2372/X U$$2505/X U$$2638/X VGND VGND VPWR VPWR dadda_fa_2_53_2/A
+ dadda_fa_2_52_5/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_45_4 U$$1693/X U$$1826/X U$$1959/X VGND VGND VPWR VPWR dadda_fa_2_46_3/B
+ dadda_fa_2_45_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_971 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_15_2 input163/X dadda_fa_4_15_2/B dadda_ha_3_15_0/SUM VGND VGND VPWR VPWR
+ dadda_fa_5_16_0/CIN dadda_fa_5_15_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1019 final_adder.U$$6/SUM final_adder.U$$505/X final_adder.U$$6/COUT
+ VGND VGND VPWR VPWR final_adder.U$$1031/B sky130_fd_sc_hd__a21o_1
XFILLER_109_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1028 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4415_1855 VGND VGND VPWR VPWR U$$4415_1855/HI U$$4415/B sky130_fd_sc_hd__conb_1
Xfanout1304 U$$3972/A VGND VGND VPWR VPWR U$$3965/B sky130_fd_sc_hd__buf_6
XFILLER_78_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1315 U$$3835/A VGND VGND VPWR VPWR U$$3828/B sky130_fd_sc_hd__buf_6
Xfanout1326 U$$955/B VGND VGND VPWR VPWR U$$958/A sky130_fd_sc_hd__buf_6
Xfanout1337 input47/X VGND VGND VPWR VPWR U$$3468/B sky130_fd_sc_hd__buf_6
Xfanout1348 U$$3425/A VGND VGND VPWR VPWR U$$3373/B sky130_fd_sc_hd__buf_6
Xfanout1359 fanout1364/X VGND VGND VPWR VPWR U$$3210/B sky130_fd_sc_hd__buf_6
XFILLER_120_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout394 U$$952/A2 VGND VGND VPWR VPWR U$$942/A2 sky130_fd_sc_hd__buf_6
XU$$3106 U$$3106/A1 U$$3108/A2 U$$3106/B1 U$$3108/B2 VGND VGND VPWR VPWR U$$3107/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3117 U$$3117/A U$$3119/B VGND VGND VPWR VPWR U$$3117/X sky130_fd_sc_hd__xor2_1
XU$$3128 U$$3948/B1 U$$3148/A2 U$$3815/A1 U$$3148/B2 VGND VGND VPWR VPWR U$$3129/A
+ sky130_fd_sc_hd__a22o_1
XU$$3139 U$$3139/A U$$3147/B VGND VGND VPWR VPWR U$$3139/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2405 U$$3775/A1 U$$2443/A2 U$$3775/B1 U$$2443/B2 VGND VGND VPWR VPWR U$$2406/A
+ sky130_fd_sc_hd__a22o_1
XU$$2416 U$$2416/A U$$2416/B VGND VGND VPWR VPWR U$$2416/X sky130_fd_sc_hd__xor2_1
XFILLER_36_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2427 U$$3112/A1 U$$2443/A2 U$$922/A1 U$$2443/B2 VGND VGND VPWR VPWR U$$2428/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2438 U$$2438/A U$$2466/A VGND VGND VPWR VPWR U$$2438/X sky130_fd_sc_hd__xor2_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2449 U$$4365/B1 U$$2459/A2 U$$4367/B1 U$$2459/B2 VGND VGND VPWR VPWR U$$2450/A
+ sky130_fd_sc_hd__a22o_1
XU$$1704 U$$882/A1 U$$1720/A2 U$$882/B1 U$$1720/B2 VGND VGND VPWR VPWR U$$1705/A sky130_fd_sc_hd__a22o_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1715 U$$1715/A U$$1721/B VGND VGND VPWR VPWR U$$1715/X sky130_fd_sc_hd__xor2_1
XU$$1726 U$$765/B1 U$$1726/A2 U$$632/A1 U$$1726/B2 VGND VGND VPWR VPWR U$$1727/A sky130_fd_sc_hd__a22o_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1737 U$$1737/A U$$1741/B VGND VGND VPWR VPWR U$$1737/X sky130_fd_sc_hd__xor2_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1748 U$$787/B1 U$$1758/A2 U$$654/A1 U$$1758/B2 VGND VGND VPWR VPWR U$$1749/A sky130_fd_sc_hd__a22o_1
XFILLER_159_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_985 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1759 U$$1759/A U$$1761/B VGND VGND VPWR VPWR U$$1759/X sky130_fd_sc_hd__xor2_1
XFILLER_15_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_316_ _321_/CLK _316_/D VGND VGND VPWR VPWR _316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput14 a[21] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__buf_4
X_247_ _247_/CLK _247_/D VGND VGND VPWR VPWR _247_/Q sky130_fd_sc_hd__dfxtp_1
Xinput25 a[31] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__buf_2
XFILLER_122_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput36 a[41] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput47 a[51] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__buf_4
XFILLER_7_864 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput58 a[61] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__clkbuf_1
X_178_ _321_/CLK _178_/D VGND VGND VPWR VPWR _178_/Q sky130_fd_sc_hd__dfxtp_1
Xinput69 b[13] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_4
XFILLER_170_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_62_4 dadda_fa_2_62_4/A dadda_fa_2_62_4/B dadda_fa_2_62_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_1/CIN dadda_fa_3_62_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_55_3 dadda_fa_2_55_3/A dadda_fa_2_55_3/B dadda_fa_2_55_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_1/B dadda_fa_3_55_3/B sky130_fd_sc_hd__fa_1
XFILLER_65_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4330 U$$4330/A U$$4350/B VGND VGND VPWR VPWR U$$4330/X sky130_fd_sc_hd__xor2_1
XU$$4341 U$$4341/A1 U$$4349/A2 U$$4480/A1 U$$4349/B2 VGND VGND VPWR VPWR U$$4342/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_48_2 dadda_fa_2_48_2/A dadda_fa_2_48_2/B dadda_fa_2_48_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_1/A dadda_fa_3_48_3/A sky130_fd_sc_hd__fa_1
XU$$4352 U$$4352/A U$$4368/B VGND VGND VPWR VPWR U$$4352/X sky130_fd_sc_hd__xor2_1
XU$$4363 U$$4363/A1 U$$4373/A2 U$$4365/A1 U$$4373/B2 VGND VGND VPWR VPWR U$$4364/A
+ sky130_fd_sc_hd__a22o_1
XU$$4374 U$$4374/A U$$4374/B VGND VGND VPWR VPWR U$$4374/X sky130_fd_sc_hd__xor2_1
XU$$4385 U$$4385/A VGND VGND VPWR VPWR U$$4387/B sky130_fd_sc_hd__inv_1
XU$$3640 U$$3775/B1 U$$3640/A2 U$$3642/A1 U$$3640/B2 VGND VGND VPWR VPWR U$$3641/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4396 U$$4396/A1 U$$4388/X U$$4398/A1 U$$4428/B2 VGND VGND VPWR VPWR U$$4397/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_25_1 dadda_fa_5_25_1/A dadda_fa_5_25_1/B dadda_fa_5_25_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_26_0/B dadda_fa_7_25_0/A sky130_fd_sc_hd__fa_1
XU$$3651 U$$3651/A U$$3695/B VGND VGND VPWR VPWR U$$3651/X sky130_fd_sc_hd__xor2_1
XU$$3662 U$$4482/B1 U$$3682/A2 U$$4349/A1 U$$3682/B2 VGND VGND VPWR VPWR U$$3663/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3673 U$$3673/A U$$3681/B VGND VGND VPWR VPWR U$$3673/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_18_0 dadda_fa_5_18_0/A dadda_fa_5_18_0/B dadda_fa_5_18_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_19_0/A dadda_fa_6_18_0/CIN sky130_fd_sc_hd__fa_1
XU$$3684 U$$3684/A1 U$$3696/A2 U$$3684/B1 U$$3696/B2 VGND VGND VPWR VPWR U$$3685/A
+ sky130_fd_sc_hd__a22o_1
XU$$3695 U$$3695/A U$$3695/B VGND VGND VPWR VPWR U$$3695/X sky130_fd_sc_hd__xor2_1
XU$$2950 U$$2950/A U$$2986/B VGND VGND VPWR VPWR U$$2950/X sky130_fd_sc_hd__xor2_1
XU$$2961 U$$3370/B1 U$$2979/A2 U$$3372/B1 U$$2979/B2 VGND VGND VPWR VPWR U$$2962/A
+ sky130_fd_sc_hd__a22o_1
XU$$2972 U$$2972/A U$$2974/B VGND VGND VPWR VPWR U$$2972/X sky130_fd_sc_hd__xor2_1
XU$$2983 U$$4353/A1 U$$3011/A2 U$$4353/B1 U$$3011/B2 VGND VGND VPWR VPWR U$$2984/A
+ sky130_fd_sc_hd__a22o_1
XU$$2994 U$$2994/A U$$3004/B VGND VGND VPWR VPWR U$$2994/X sky130_fd_sc_hd__xor2_1
XFILLER_138_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$901 final_adder.U$$130/A final_adder.U$$839/X final_adder.U$$901/B1
+ VGND VGND VPWR VPWR final_adder.U$$901/X sky130_fd_sc_hd__a21o_1
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$923 final_adder.U$$152/A final_adder.U$$861/X final_adder.U$$923/B1
+ VGND VGND VPWR VPWR final_adder.U$$923/X sky130_fd_sc_hd__a21o_1
XFILLER_113_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$945 final_adder.U$$174/A final_adder.U$$883/X final_adder.U$$945/B1
+ VGND VGND VPWR VPWR final_adder.U$$945/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_2 U$$905/X U$$1038/X U$$1171/X VGND VGND VPWR VPWR dadda_fa_2_51_1/A
+ dadda_fa_2_50_4/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$967 final_adder.U$$196/A final_adder.U$$809/X final_adder.U$$967/B1
+ VGND VGND VPWR VPWR final_adder.U$$967/X sky130_fd_sc_hd__a21o_1
XU$$806 U$$806/A U$$822/A VGND VGND VPWR VPWR U$$806/X sky130_fd_sc_hd__xor2_1
XU$$817 U$$954/A1 U$$817/A2 U$$956/A1 U$$817/B2 VGND VGND VPWR VPWR U$$818/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_43_1 U$$492/X U$$625/X U$$758/X VGND VGND VPWR VPWR dadda_fa_2_44_3/A
+ dadda_fa_2_43_5/A sky130_fd_sc_hd__fa_1
XFILLER_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$989 final_adder.U$$218/A final_adder.U$$831/X final_adder.U$$989/B1
+ VGND VGND VPWR VPWR final_adder.U$$989/X sky130_fd_sc_hd__a21o_1
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$828 U$$828/A1 U$$910/A2 U$$828/B1 U$$910/B2 VGND VGND VPWR VPWR U$$829/A sky130_fd_sc_hd__a22o_1
XFILLER_83_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$839 U$$839/A U$$907/B VGND VGND VPWR VPWR U$$839/X sky130_fd_sc_hd__xor2_1
XFILLER_16_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_20_0 U$$1449/B input169/X dadda_fa_4_20_0/CIN VGND VGND VPWR VPWR dadda_fa_5_21_0/A
+ dadda_fa_5_20_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_36_0 U$$79/X U$$212/X U$$345/X VGND VGND VPWR VPWR dadda_fa_2_37_5/A dadda_fa_2_36_5/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_169_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_72_3 dadda_fa_3_72_3/A dadda_fa_3_72_3/B dadda_fa_3_72_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_1/B dadda_fa_4_72_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1101 input81/X VGND VGND VPWR VPWR U$$3618/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_65_2 dadda_fa_3_65_2/A dadda_fa_3_65_2/B dadda_fa_3_65_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_1/A dadda_fa_4_65_2/B sky130_fd_sc_hd__fa_1
Xfanout1112 input79/X VGND VGND VPWR VPWR U$$735/B1 sky130_fd_sc_hd__buf_4
Xfanout1123 U$$4434/A1 VGND VGND VPWR VPWR U$$4295/B1 sky130_fd_sc_hd__buf_6
Xfanout1134 U$$3296/B1 VGND VGND VPWR VPWR U$$3022/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1145 input75/X VGND VGND VPWR VPWR U$$4430/A1 sky130_fd_sc_hd__buf_4
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1156 U$$316/B1 VGND VGND VPWR VPWR U$$2647/A1 sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_3_58_1 dadda_fa_3_58_1/A dadda_fa_3_58_1/B dadda_fa_3_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_0/CIN dadda_fa_4_58_2/A sky130_fd_sc_hd__fa_1
Xfanout1167 input73/X VGND VGND VPWR VPWR U$$4424/B1 sky130_fd_sc_hd__buf_4
XFILLER_120_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1178 U$$3189/A1 VGND VGND VPWR VPWR U$$721/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_6_35_0 dadda_fa_6_35_0/A dadda_fa_6_35_0/B dadda_fa_6_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_36_0/B dadda_fa_7_35_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1189 U$$3048/B1 VGND VGND VPWR VPWR U$$36/A1 sky130_fd_sc_hd__buf_4
XFILLER_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2202 U$$969/A1 U$$2252/A2 U$$971/A1 U$$2252/B2 VGND VGND VPWR VPWR U$$2203/A sky130_fd_sc_hd__a22o_1
XFILLER_62_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2213 U$$2213/A U$$2253/B VGND VGND VPWR VPWR U$$2213/X sky130_fd_sc_hd__xor2_1
XU$$2224 U$$991/A1 U$$2254/A2 U$$993/A1 U$$2254/B2 VGND VGND VPWR VPWR U$$2225/A sky130_fd_sc_hd__a22o_1
XU$$2235 U$$2235/A U$$2253/B VGND VGND VPWR VPWR U$$2235/X sky130_fd_sc_hd__xor2_1
XU$$1501 U$$1501/A U$$1507/A VGND VGND VPWR VPWR U$$1501/X sky130_fd_sc_hd__xor2_1
XFILLER_16_941 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2246 U$$739/A1 U$$2248/A2 U$$741/A1 U$$2248/B2 VGND VGND VPWR VPWR U$$2247/A sky130_fd_sc_hd__a22o_1
XU$$1512 U$$1510/B U$$1497/B input15/X U$$1507/Y VGND VGND VPWR VPWR U$$1512/X sky130_fd_sc_hd__a22o_1
XFILLER_62_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2257 U$$2257/A U$$2269/B VGND VGND VPWR VPWR U$$2257/X sky130_fd_sc_hd__xor2_1
XFILLER_34_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1523 U$$2891/B1 U$$1563/A2 U$$2758/A1 U$$1563/B2 VGND VGND VPWR VPWR U$$1524/A
+ sky130_fd_sc_hd__a22o_1
XU$$2268 U$$487/A1 U$$2272/A2 U$$487/B1 U$$2272/B2 VGND VGND VPWR VPWR U$$2269/A sky130_fd_sc_hd__a22o_1
XU$$1534 U$$1534/A U$$1570/B VGND VGND VPWR VPWR U$$1534/X sky130_fd_sc_hd__xor2_1
XU$$2279 U$$2279/A U$$2283/B VGND VGND VPWR VPWR U$$2279/X sky130_fd_sc_hd__xor2_1
XU$$1545 U$$38/A1 U$$1575/A2 U$$40/A1 U$$1575/B2 VGND VGND VPWR VPWR U$$1546/A sky130_fd_sc_hd__a22o_1
XU$$1556 U$$1556/A U$$1564/B VGND VGND VPWR VPWR U$$1556/X sky130_fd_sc_hd__xor2_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1567 U$$469/B1 U$$1567/A2 U$$884/A1 U$$1567/B2 VGND VGND VPWR VPWR U$$1568/A sky130_fd_sc_hd__a22o_1
XFILLER_31_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1578 U$$1578/A U$$1584/B VGND VGND VPWR VPWR U$$1578/X sky130_fd_sc_hd__xor2_1
XU$$1589 U$$765/B1 U$$1593/A2 U$$632/A1 U$$1593/B2 VGND VGND VPWR VPWR U$$1590/A sky130_fd_sc_hd__a22o_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_108_0 dadda_fa_7_108_0/A dadda_fa_7_108_0/B dadda_fa_7_108_0/CIN VGND
+ VGND VPWR VPWR _405_/D _276_/D sky130_fd_sc_hd__fa_1
XFILLER_156_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_1 dadda_fa_2_60_1/A dadda_fa_2_60_1/B dadda_fa_2_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_0/CIN dadda_fa_3_60_2/CIN sky130_fd_sc_hd__fa_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$208 final_adder.U$$208/A final_adder.U$$208/B VGND VGND VPWR VPWR
+ final_adder.U$$336/B sky130_fd_sc_hd__and2_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$219 final_adder.U$$218/B final_adder.U$$989/B1 final_adder.U$$219/B1
+ VGND VGND VPWR VPWR final_adder.U$$219/X sky130_fd_sc_hd__a21o_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_53_0 dadda_fa_2_53_0/A dadda_fa_2_53_0/B dadda_fa_2_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_0/B dadda_fa_3_53_2/B sky130_fd_sc_hd__fa_1
Xfanout1690 U$$1360/B VGND VGND VPWR VPWR U$$1358/B sky130_fd_sc_hd__buf_8
XU$$4160 U$$4295/B1 U$$4174/A2 U$$4162/A1 U$$4174/B2 VGND VGND VPWR VPWR U$$4161/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4171 U$$4171/A U$$4175/B VGND VGND VPWR VPWR U$$4171/X sky130_fd_sc_hd__xor2_1
XFILLER_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4182 U$$4182/A1 U$$4240/A2 U$$4458/A1 U$$4240/B2 VGND VGND VPWR VPWR U$$4183/A
+ sky130_fd_sc_hd__a22o_1
XU$$4193 U$$4193/A U$$4215/B VGND VGND VPWR VPWR U$$4193/X sky130_fd_sc_hd__xor2_1
XU$$3470 U$$3470/A U$$3474/B VGND VGND VPWR VPWR U$$3470/X sky130_fd_sc_hd__xor2_1
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3481 U$$3618/A1 U$$3523/A2 U$$3618/B1 U$$3523/B2 VGND VGND VPWR VPWR U$$3482/A
+ sky130_fd_sc_hd__a22o_1
XU$$3492 U$$3492/A U$$3506/B VGND VGND VPWR VPWR U$$3492/X sky130_fd_sc_hd__xor2_1
XFILLER_41_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2780 U$$2780/A1 U$$2856/A2 U$$2780/B1 U$$2856/B2 VGND VGND VPWR VPWR U$$2781/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_7_0 U$$21/X U$$154/X U$$287/X VGND VGND VPWR VPWR dadda_fa_6_8_0/A dadda_fa_6_7_0/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_22_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2791 U$$2791/A U$$2799/B VGND VGND VPWR VPWR U$$2791/X sky130_fd_sc_hd__xor2_1
XFILLER_139_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_82_2 dadda_fa_4_82_2/A dadda_fa_4_82_2/B dadda_fa_4_82_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_83_0/CIN dadda_fa_5_82_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_75_1 dadda_fa_4_75_1/A dadda_fa_4_75_1/B dadda_fa_4_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_76_0/B dadda_fa_5_75_1/B sky130_fd_sc_hd__fa_1
XFILLER_161_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_52_0 dadda_fa_7_52_0/A dadda_fa_7_52_0/B dadda_fa_7_52_0/CIN VGND VGND
+ VPWR VPWR _349_/D _220_/D sky130_fd_sc_hd__fa_1
XFILLER_161_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_68_0 dadda_fa_4_68_0/A dadda_fa_4_68_0/B dadda_fa_4_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_69_0/A dadda_fa_5_68_1/A sky130_fd_sc_hd__fa_1
Xinput204 c[52] VGND VGND VPWR VPWR input204/X sky130_fd_sc_hd__buf_2
XFILLER_89_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput215 c[62] VGND VGND VPWR VPWR input215/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput226 c[72] VGND VGND VPWR VPWR input226/X sky130_fd_sc_hd__buf_2
Xinput237 c[82] VGND VGND VPWR VPWR input237/X sky130_fd_sc_hd__clkbuf_1
Xinput248 c[92] VGND VGND VPWR VPWR input248/X sky130_fd_sc_hd__buf_2
XFILLER_25_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$720 final_adder.U$$720/A final_adder.U$$720/B VGND VGND VPWR VPWR
+ final_adder.U$$800/A sky130_fd_sc_hd__and2_1
XFILLER_29_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$731 final_adder.U$$714/A final_adder.U$$503/X final_adder.U$$611/X
+ VGND VGND VPWR VPWR final_adder.U$$731/X sky130_fd_sc_hd__a21o_2
XFILLER_57_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$742 final_adder.U$$774/B final_adder.U$$742/B VGND VGND VPWR VPWR
+ final_adder.U$$742/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$753 final_adder.U$$752/B final_adder.U$$673/X final_adder.U$$641/X
+ VGND VGND VPWR VPWR final_adder.U$$753/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$764 final_adder.U$$796/B final_adder.U$$764/B VGND VGND VPWR VPWR
+ final_adder.U$$764/X sky130_fd_sc_hd__and2_1
XFILLER_56_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$603 U$$603/A U$$637/B VGND VGND VPWR VPWR U$$603/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$775 final_adder.U$$774/B final_adder.U$$695/X final_adder.U$$663/X
+ VGND VGND VPWR VPWR final_adder.U$$775/X sky130_fd_sc_hd__a21o_1
XU$$614 U$$749/B1 U$$638/A2 U$$616/A1 U$$638/B2 VGND VGND VPWR VPWR U$$615/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$786 final_adder.U$$786/A final_adder.U$$786/B VGND VGND VPWR VPWR
+ final_adder.U$$786/X sky130_fd_sc_hd__and2_1
XU$$625 U$$625/A U$$631/B VGND VGND VPWR VPWR U$$625/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$797 final_adder.U$$796/B final_adder.U$$717/X final_adder.U$$685/X
+ VGND VGND VPWR VPWR final_adder.U$$797/X sky130_fd_sc_hd__a21o_1
XU$$636 U$$88/A1 U$$636/A2 U$$88/B1 U$$636/B2 VGND VGND VPWR VPWR U$$637/A sky130_fd_sc_hd__a22o_1
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$647 U$$647/A U$$684/A VGND VGND VPWR VPWR U$$647/X sky130_fd_sc_hd__xor2_1
XU$$658 U$$932/A1 U$$674/A2 U$$934/A1 U$$674/B2 VGND VGND VPWR VPWR U$$659/A sky130_fd_sc_hd__a22o_1
XFILLER_83_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$669 U$$669/A U$$669/B VGND VGND VPWR VPWR U$$669/X sky130_fd_sc_hd__xor2_1
XFILLER_71_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_70_0 dadda_fa_3_70_0/A dadda_fa_3_70_0/B dadda_fa_3_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_0/B dadda_fa_4_70_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2010 U$$640/A1 U$$2052/A2 U$$916/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2011/A sky130_fd_sc_hd__a22o_1
XU$$4467_1881 VGND VGND VPWR VPWR U$$4467_1881/HI U$$4467/B sky130_fd_sc_hd__conb_1
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2021 U$$2021/A U$$2053/B VGND VGND VPWR VPWR U$$2021/X sky130_fd_sc_hd__xor2_1
XU$$2032 U$$388/A1 U$$2046/A2 U$$2443/B1 U$$2046/B2 VGND VGND VPWR VPWR U$$2033/A
+ sky130_fd_sc_hd__a22o_1
XU$$2043 U$$2043/A U$$2043/B VGND VGND VPWR VPWR U$$2043/X sky130_fd_sc_hd__xor2_1
XU$$2054 U$$2054/A VGND VGND VPWR VPWR U$$2054/Y sky130_fd_sc_hd__inv_1
XFILLER_50_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2065 U$$3296/B1 U$$2097/A2 U$$3298/B1 U$$2097/B2 VGND VGND VPWR VPWR U$$2066/A
+ sky130_fd_sc_hd__a22o_1
XU$$1320 U$$1320/A U$$1320/B VGND VGND VPWR VPWR U$$1320/X sky130_fd_sc_hd__xor2_1
XU$$1331 U$$2973/B1 U$$1367/A2 U$$98/B1 U$$1367/B2 VGND VGND VPWR VPWR U$$1332/A sky130_fd_sc_hd__a22o_1
XU$$2076 U$$2076/A U$$2106/B VGND VGND VPWR VPWR U$$2076/X sky130_fd_sc_hd__xor2_1
XU$$2087 U$$991/A1 U$$2097/A2 U$$993/A1 U$$2097/B2 VGND VGND VPWR VPWR U$$2088/A sky130_fd_sc_hd__a22o_1
XU$$1342 U$$1342/A U$$1364/B VGND VGND VPWR VPWR U$$1342/X sky130_fd_sc_hd__xor2_1
XFILLER_16_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2098 U$$2098/A U$$2130/B VGND VGND VPWR VPWR U$$2098/X sky130_fd_sc_hd__xor2_1
XU$$1353 U$$120/A1 U$$1353/A2 U$$120/B1 U$$1353/B2 VGND VGND VPWR VPWR U$$1354/A sky130_fd_sc_hd__a22o_1
XU$$1364 U$$1364/A U$$1364/B VGND VGND VPWR VPWR U$$1364/X sky130_fd_sc_hd__xor2_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1375 U$$1373/B U$$1370/A input13/X U$$1370/Y VGND VGND VPWR VPWR U$$1375/X sky130_fd_sc_hd__a22o_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_916 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1386 U$$3030/A1 U$$1432/A2 U$$3030/B1 U$$1432/B2 VGND VGND VPWR VPWR U$$1387/A
+ sky130_fd_sc_hd__a22o_1
XU$$1397 U$$1397/A U$$1433/B VGND VGND VPWR VPWR U$$1397/X sky130_fd_sc_hd__xor2_1
XFILLER_157_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_92_1 dadda_fa_5_92_1/A dadda_fa_5_92_1/B dadda_fa_5_92_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_93_0/B dadda_fa_7_92_0/A sky130_fd_sc_hd__fa_1
XFILLER_159_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_85_0 dadda_fa_5_85_0/A dadda_fa_5_85_0/B dadda_fa_5_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_86_0/A dadda_fa_6_85_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_104_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout905 U$$1202/B2 VGND VGND VPWR VPWR U$$1194/B2 sky130_fd_sc_hd__buf_4
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout916 U$$80/B2 VGND VGND VPWR VPWR U$$48/B2 sky130_fd_sc_hd__buf_2
Xfanout927 U$$4502/B2 VGND VGND VPWR VPWR U$$4492/B2 sky130_fd_sc_hd__buf_2
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_77_7 U$$4151/X U$$4284/X U$$4417/X VGND VGND VPWR VPWR dadda_fa_2_78_2/CIN
+ dadda_fa_2_77_5/CIN sky130_fd_sc_hd__fa_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout938 input99/X VGND VGND VPWR VPWR fanout938/X sky130_fd_sc_hd__buf_6
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout949 fanout957/X VGND VGND VPWR VPWR U$$632/B1 sky130_fd_sc_hd__buf_4
XFILLER_86_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$60 _356_/Q _228_/Q VGND VGND VPWR VPWR final_adder.U$$965/B1 final_adder.U$$194/A
+ sky130_fd_sc_hd__ha_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$71 _367_/Q _239_/Q VGND VGND VPWR VPWR final_adder.U$$185/B1 final_adder.U$$184/B
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$82 _378_/Q _250_/Q VGND VGND VPWR VPWR final_adder.U$$943/B1 final_adder.U$$172/A
+ sky130_fd_sc_hd__ha_1
XFILLER_53_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$93 _389_/Q _261_/Q VGND VGND VPWR VPWR final_adder.U$$163/B1 final_adder.U$$162/B
+ sky130_fd_sc_hd__ha_1
XFILLER_13_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_101_2 dadda_fa_3_101_2/A dadda_fa_3_101_2/B dadda_fa_3_101_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_102_1/A dadda_fa_4_101_2/B sky130_fd_sc_hd__fa_1
XFILLER_79_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_65_5 U$$2132/X U$$2265/X U$$2398/X VGND VGND VPWR VPWR dadda_fa_1_66_7/A
+ dadda_fa_2_65_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_115_0 dadda_fa_6_115_0/A dadda_fa_6_115_0/B dadda_fa_6_115_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_116_0/B dadda_fa_7_115_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$550 final_adder.U$$558/B final_adder.U$$550/B VGND VGND VPWR VPWR
+ final_adder.U$$670/B sky130_fd_sc_hd__and2_1
XFILLER_57_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$561 final_adder.U$$560/B final_adder.U$$445/X final_adder.U$$437/X
+ VGND VGND VPWR VPWR final_adder.U$$561/X sky130_fd_sc_hd__a21o_1
XU$$400 U$$672/B1 U$$406/A2 U$$539/A1 U$$406/B2 VGND VGND VPWR VPWR U$$401/A sky130_fd_sc_hd__a22o_1
XFILLER_85_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$572 final_adder.U$$580/B final_adder.U$$572/B VGND VGND VPWR VPWR
+ final_adder.U$$692/B sky130_fd_sc_hd__and2_1
XU$$411 U$$411/A VGND VGND VPWR VPWR U$$411/Y sky130_fd_sc_hd__inv_1
XFILLER_63_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$583 final_adder.U$$582/B final_adder.U$$467/X final_adder.U$$459/X
+ VGND VGND VPWR VPWR final_adder.U$$583/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_3_35_3 dadda_fa_3_35_3/A dadda_fa_3_35_3/B dadda_fa_3_35_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_1/B dadda_fa_4_35_2/CIN sky130_fd_sc_hd__fa_1
XU$$422 U$$422/A U$$448/B VGND VGND VPWR VPWR U$$422/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$594 final_adder.U$$602/B final_adder.U$$594/B VGND VGND VPWR VPWR
+ final_adder.U$$714/B sky130_fd_sc_hd__and2_1
XU$$433 U$$22/A1 U$$447/A2 U$$24/A1 U$$447/B2 VGND VGND VPWR VPWR U$$434/A sky130_fd_sc_hd__a22o_1
XU$$444 U$$444/A U$$506/B VGND VGND VPWR VPWR U$$444/X sky130_fd_sc_hd__xor2_1
XU$$455 U$$864/B1 U$$497/A2 U$$729/B1 U$$497/B2 VGND VGND VPWR VPWR U$$456/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_28_2 dadda_fa_3_28_2/A dadda_fa_3_28_2/B dadda_fa_3_28_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_29_1/A dadda_fa_4_28_2/B sky130_fd_sc_hd__fa_1
XFILLER_45_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$466 U$$466/A U$$504/B VGND VGND VPWR VPWR U$$466/X sky130_fd_sc_hd__xor2_1
XFILLER_72_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$477 U$$612/B1 U$$479/A2 U$$479/A1 U$$479/B2 VGND VGND VPWR VPWR U$$478/A sky130_fd_sc_hd__a22o_1
XU$$488 U$$488/A U$$504/B VGND VGND VPWR VPWR U$$488/X sky130_fd_sc_hd__xor2_1
XFILLER_60_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$499 U$$499/A1 U$$539/A2 U$$90/A1 U$$539/B2 VGND VGND VPWR VPWR U$$500/A sky130_fd_sc_hd__a22o_1
XFILLER_60_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4497_1896 VGND VGND VPWR VPWR U$$4497_1896/HI U$$4497/B sky130_fd_sc_hd__conb_1
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_2_31_4 U$$1665/X U$$1798/X VGND VGND VPWR VPWR dadda_fa_3_32_2/A dadda_fa_4_31_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_121_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_7_1_0 U$$9/X input168/X VGND VGND VPWR VPWR _298_/D _169_/D sky130_fd_sc_hd__ha_1
XFILLER_94_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_30_2 U$$865/X U$$998/X U$$1131/X VGND VGND VPWR VPWR dadda_fa_3_31_1/CIN
+ dadda_fa_3_30_3/B sky130_fd_sc_hd__fa_2
XFILLER_36_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1150 U$$54/A1 U$$1194/A2 U$$56/A1 U$$1194/B2 VGND VGND VPWR VPWR U$$1151/A sky130_fd_sc_hd__a22o_1
XU$$1161 U$$1161/A U$$1163/B VGND VGND VPWR VPWR U$$1161/X sky130_fd_sc_hd__xor2_1
XU$$1172 U$$74/B1 U$$1174/A2 U$$215/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1173/A sky130_fd_sc_hd__a22o_1
XU$$1183 U$$1183/A U$$1227/B VGND VGND VPWR VPWR U$$1183/X sky130_fd_sc_hd__xor2_1
XU$$1194 U$$98/A1 U$$1194/A2 U$$98/B1 U$$1194/B2 VGND VGND VPWR VPWR U$$1195/A sky130_fd_sc_hd__a22o_1
XU$$2326_1801 VGND VGND VPWR VPWR U$$2326_1801/HI U$$2326/B1 sky130_fd_sc_hd__conb_1
XFILLER_136_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_82_5 U$$3230/X U$$3363/X U$$3496/X VGND VGND VPWR VPWR dadda_fa_2_83_3/A
+ dadda_fa_2_82_5/B sky130_fd_sc_hd__fa_1
Xfanout702 U$$4244/B2 VGND VGND VPWR VPWR U$$4174/B2 sky130_fd_sc_hd__buf_4
Xfanout713 U$$4057/B2 VGND VGND VPWR VPWR U$$4105/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_172_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_75_4 U$$3216/X U$$3349/X U$$3482/X VGND VGND VPWR VPWR dadda_fa_2_76_1/CIN
+ dadda_fa_2_75_4/CIN sky130_fd_sc_hd__fa_1
Xfanout724 U$$3966/B2 VGND VGND VPWR VPWR U$$3960/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout735 U$$3644/B2 VGND VGND VPWR VPWR U$$3604/B2 sky130_fd_sc_hd__buf_4
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout746 U$$3430/X VGND VGND VPWR VPWR U$$3473/B2 sky130_fd_sc_hd__buf_4
XFILLER_113_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout757 U$$3422/B2 VGND VGND VPWR VPWR U$$3416/B2 sky130_fd_sc_hd__buf_4
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_3 U$$3734/X U$$3867/X U$$4000/X VGND VGND VPWR VPWR dadda_fa_2_69_1/B
+ dadda_fa_2_68_4/B sky130_fd_sc_hd__fa_1
Xfanout768 U$$3257/B2 VGND VGND VPWR VPWR U$$3251/B2 sky130_fd_sc_hd__buf_2
XFILLER_100_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout779 U$$2937/B2 VGND VGND VPWR VPWR U$$2929/B2 sky130_fd_sc_hd__buf_4
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_45_2 dadda_fa_4_45_2/A dadda_fa_4_45_2/B dadda_fa_4_45_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_46_0/CIN dadda_fa_5_45_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_38_1 dadda_fa_4_38_1/A dadda_fa_4_38_1/B dadda_fa_4_38_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_39_0/B dadda_fa_5_38_1/B sky130_fd_sc_hd__fa_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_15_0 dadda_fa_7_15_0/A dadda_fa_7_15_0/B dadda_fa_7_15_0/CIN VGND VGND
+ VPWR VPWR _312_/D _183_/D sky130_fd_sc_hd__fa_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_280_ _416_/CLK _280_/D VGND VGND VPWR VPWR _280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_70_3 U$$1610/X U$$1743/X U$$1876/X VGND VGND VPWR VPWR dadda_fa_1_71_7/B
+ dadda_fa_1_70_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_7_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_63_2 U$$931/X U$$1064/X U$$1197/X VGND VGND VPWR VPWR dadda_fa_1_64_6/A
+ dadda_fa_1_63_8/A sky130_fd_sc_hd__fa_1
XFILLER_37_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_40_1 dadda_fa_3_40_1/A dadda_fa_3_40_1/B dadda_fa_3_40_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_0/CIN dadda_fa_4_40_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_0_56_1 U$$518/X U$$651/X U$$784/X VGND VGND VPWR VPWR dadda_fa_1_57_7/CIN
+ dadda_fa_1_56_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_64_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_33_0 input183/X dadda_fa_3_33_0/B dadda_fa_3_33_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_34_0/B dadda_fa_4_33_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_92_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$230 U$$230/A U$$230/B VGND VGND VPWR VPWR U$$230/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$391 final_adder.U$$390/B final_adder.U$$269/X final_adder.U$$265/X
+ VGND VGND VPWR VPWR final_adder.U$$391/X sky130_fd_sc_hd__a21o_1
XU$$241 U$$787/B1 U$$253/A2 U$$654/A1 U$$253/B2 VGND VGND VPWR VPWR U$$242/A sky130_fd_sc_hd__a22o_1
XU$$252 U$$252/A U$$254/B VGND VGND VPWR VPWR U$$252/X sky130_fd_sc_hd__xor2_1
XU$$263 U$$672/B1 U$$271/A2 U$$539/A1 U$$271/B2 VGND VGND VPWR VPWR U$$264/A sky130_fd_sc_hd__a22o_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$274 U$$274/A VGND VGND VPWR VPWR U$$274/Y sky130_fd_sc_hd__inv_1
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$285 U$$285/A U$$313/B VGND VGND VPWR VPWR U$$285/X sky130_fd_sc_hd__xor2_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$296 U$$22/A1 U$$312/A2 U$$24/A1 U$$312/B2 VGND VGND VPWR VPWR U$$297/A sky130_fd_sc_hd__a22o_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2 U$$3/A VGND VGND VPWR VPWR U$$2/Y sky130_fd_sc_hd__inv_1
XFILLER_69_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput305 output305/A VGND VGND VPWR VPWR o[28] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_4 input248/X dadda_fa_2_92_4/B dadda_fa_2_92_4/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_93_1/CIN dadda_fa_3_92_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput316 output316/A VGND VGND VPWR VPWR o[38] sky130_fd_sc_hd__buf_2
Xoutput327 output327/A VGND VGND VPWR VPWR o[48] sky130_fd_sc_hd__buf_2
Xoutput338 output338/A VGND VGND VPWR VPWR o[58] sky130_fd_sc_hd__buf_2
Xoutput349 output349/A VGND VGND VPWR VPWR o[68] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_85_3 dadda_fa_2_85_3/A dadda_fa_2_85_3/B dadda_fa_2_85_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_1/B dadda_fa_3_85_3/B sky130_fd_sc_hd__fa_1
XFILLER_126_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_78_2 dadda_fa_2_78_2/A dadda_fa_2_78_2/B dadda_fa_2_78_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_1/A dadda_fa_3_78_3/A sky130_fd_sc_hd__fa_1
XFILLER_141_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_55_1 dadda_fa_5_55_1/A dadda_fa_5_55_1/B dadda_fa_5_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_56_0/B dadda_fa_7_55_0/A sky130_fd_sc_hd__fa_1
XFILLER_141_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_48_0 dadda_fa_5_48_0/A dadda_fa_5_48_0/B dadda_fa_5_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_49_0/A dadda_fa_6_48_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_ha_2_22_0 U$$51/X U$$184/X VGND VGND VPWR VPWR dadda_fa_3_23_3/CIN dadda_fa_4_22_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_132_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_47_clk _218_/CLK VGND VGND VPWR VPWR _348_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_101_1 U$$3002/X U$$3135/X U$$3268/X VGND VGND VPWR VPWR dadda_fa_3_102_2/A
+ dadda_fa_3_101_3/B sky130_fd_sc_hd__fa_1
XFILLER_50_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_122_0 U$$4241/X U$$4374/X U$$4507/X VGND VGND VPWR VPWR dadda_fa_6_123_0/A
+ dadda_fa_6_122_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_80_2 U$$1896/X U$$2029/X U$$2162/X VGND VGND VPWR VPWR dadda_fa_2_81_1/B
+ dadda_fa_2_80_4/A sky130_fd_sc_hd__fa_1
XFILLER_120_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout510 U$$3155/X VGND VGND VPWR VPWR U$$3257/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout1508 U$$985/A1 VGND VGND VPWR VPWR U$$3999/A1 sky130_fd_sc_hd__buf_4
Xfanout521 U$$2977/A2 VGND VGND VPWR VPWR U$$2937/A2 sky130_fd_sc_hd__buf_6
Xfanout1519 U$$3447/B1 VGND VGND VPWR VPWR U$$709/A1 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_1_73_1 U$$2281/X U$$2414/X U$$2547/X VGND VGND VPWR VPWR dadda_fa_2_74_0/CIN
+ dadda_fa_2_73_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout532 U$$340/A2 VGND VGND VPWR VPWR U$$312/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout543 U$$2812/A2 VGND VGND VPWR VPWR U$$2874/A2 sky130_fd_sc_hd__buf_6
Xfanout554 fanout561/X VGND VGND VPWR VPWR U$$2540/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_4_50_0 dadda_fa_4_50_0/A dadda_fa_4_50_0/B dadda_fa_4_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_51_0/A dadda_fa_5_50_1/A sky130_fd_sc_hd__fa_1
XFILLER_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout565 U$$2333/X VGND VGND VPWR VPWR U$$2445/A2 sky130_fd_sc_hd__buf_4
XFILLER_101_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_66_0 U$$2533/X U$$2666/X U$$2799/X VGND VGND VPWR VPWR dadda_fa_2_67_0/B
+ dadda_fa_2_66_3/B sky130_fd_sc_hd__fa_1
XFILLER_76_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout576 U$$2320/A2 VGND VGND VPWR VPWR U$$2326/A2 sky130_fd_sc_hd__clkbuf_8
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout587 U$$2014/A2 VGND VGND VPWR VPWR U$$1986/A2 sky130_fd_sc_hd__buf_4
Xfanout598 U$$1891/A2 VGND VGND VPWR VPWR U$$1881/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_100_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_38_clk _388_/CLK VGND VGND VPWR VPWR _369_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$2609 U$$2609/A1 U$$2681/A2 U$$967/A1 U$$2681/B2 VGND VGND VPWR VPWR U$$2610/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1908 U$$1908/A U$$1910/B VGND VGND VPWR VPWR U$$1908/X sky130_fd_sc_hd__xor2_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_401_ _402_/CLK _401_/D VGND VGND VPWR VPWR _401_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1919 input21/X VGND VGND VPWR VPWR U$$1921/B sky130_fd_sc_hd__inv_1
XFILLER_42_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_332_ _344_/CLK _332_/D VGND VGND VPWR VPWR _332_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_263_ _391_/CLK _263_/D VGND VGND VPWR VPWR _263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_194_ _328_/CLK _194_/D VGND VGND VPWR VPWR _194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_95_2 dadda_fa_3_95_2/A dadda_fa_3_95_2/B dadda_fa_3_95_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_1/A dadda_fa_4_95_2/B sky130_fd_sc_hd__fa_1
XFILLER_109_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_88_1 dadda_fa_3_88_1/A dadda_fa_3_88_1/B dadda_fa_3_88_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_0/CIN dadda_fa_4_88_2/A sky130_fd_sc_hd__fa_1
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_65_0 dadda_fa_6_65_0/A dadda_fa_6_65_0/B dadda_fa_6_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_66_0/B dadda_fa_7_65_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_44_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4390_1842 VGND VGND VPWR VPWR U$$4390_1842/HI U$$4390/A1 sky130_fd_sc_hd__conb_1
XFILLER_97_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4501 U$$4501/A U$$4501/B VGND VGND VPWR VPWR U$$4501/X sky130_fd_sc_hd__xor2_1
XFILLER_65_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4512 U$$4512/A1 U$$4388/X U$$4512/B1 U$$4516/B2 VGND VGND VPWR VPWR U$$4513/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3800 U$$3800/A U$$3816/B VGND VGND VPWR VPWR U$$3800/X sky130_fd_sc_hd__xor2_1
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$15 U$$15/A U$$9/B VGND VGND VPWR VPWR U$$15/X sky130_fd_sc_hd__xor2_1
XFILLER_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3811 U$$3948/A1 U$$3825/A2 U$$3948/B1 U$$3825/B2 VGND VGND VPWR VPWR U$$3812/A
+ sky130_fd_sc_hd__a22o_1
XU$$26 U$$26/A1 U$$48/A2 U$$28/A1 U$$48/B2 VGND VGND VPWR VPWR U$$27/A sky130_fd_sc_hd__a22o_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$37 U$$37/A U$$77/B VGND VGND VPWR VPWR U$$37/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_117_1 U$$4098/X U$$4231/X U$$4364/X VGND VGND VPWR VPWR dadda_fa_5_118_0/B
+ dadda_fa_5_117_1/B sky130_fd_sc_hd__fa_1
XU$$3822 U$$3822/A U$$3828/B VGND VGND VPWR VPWR U$$3822/X sky130_fd_sc_hd__xor2_1
XFILLER_53_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3833 U$$3833/A1 U$$3833/A2 U$$3833/B1 U$$3833/B2 VGND VGND VPWR VPWR U$$3834/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3844 U$$3979/B1 U$$3924/A2 U$$3846/A1 U$$3924/B2 VGND VGND VPWR VPWR U$$3845/A
+ sky130_fd_sc_hd__a22o_1
XU$$48 U$$48/A1 U$$48/A2 U$$50/A1 U$$48/B2 VGND VGND VPWR VPWR U$$49/A sky130_fd_sc_hd__a22o_1
XU$$3855 U$$3855/A U$$3867/B VGND VGND VPWR VPWR U$$3855/X sky130_fd_sc_hd__xor2_1
XU$$59 U$$59/A U$$97/B VGND VGND VPWR VPWR U$$59/X sky130_fd_sc_hd__xor2_1
XFILLER_46_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3866 U$$4001/B1 U$$3892/A2 U$$854/A1 U$$3892/B2 VGND VGND VPWR VPWR U$$3867/A
+ sky130_fd_sc_hd__a22o_1
XU$$3877 U$$3877/A U$$3925/B VGND VGND VPWR VPWR U$$3877/X sky130_fd_sc_hd__xor2_1
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3888 U$$4162/A1 U$$3906/A2 U$$4162/B1 U$$3906/B2 VGND VGND VPWR VPWR U$$3889/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3899 U$$3899/A U$$3907/B VGND VGND VPWR VPWR U$$3899/X sky130_fd_sc_hd__xor2_1
XFILLER_61_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_90_1 U$$3645/X U$$3778/X U$$3911/X VGND VGND VPWR VPWR dadda_fa_3_91_0/CIN
+ dadda_fa_3_90_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_83_0 U$$4163/X U$$4296/X U$$4429/X VGND VGND VPWR VPWR dadda_fa_3_84_0/B
+ dadda_fa_3_83_2/B sky130_fd_sc_hd__fa_1
XFILLER_102_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_52_6 U$$2771/X U$$2904/X U$$3037/X VGND VGND VPWR VPWR dadda_fa_2_53_2/B
+ dadda_fa_2_52_5/B sky130_fd_sc_hd__fa_1
XFILLER_56_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_983 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_4_0 dadda_fa_7_4_0/A dadda_fa_7_4_0/B dadda_fa_7_4_0/CIN VGND VGND VPWR
+ VPWR _301_/D _172_/D sky130_fd_sc_hd__fa_1
XFILLER_36_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_5_126_0_1947 VGND VGND VPWR VPWR dadda_ha_5_126_0/A dadda_ha_5_126_0_1947/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1009 final_adder.U$$238/A final_adder.U$$619/X final_adder.U$$239/A2
+ VGND VGND VPWR VPWR final_adder.U$$1041/B sky130_fd_sc_hd__a21o_1
XFILLER_137_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_82_0 dadda_fa_7_82_0/A dadda_fa_7_82_0/B dadda_fa_7_82_0/CIN VGND VGND
+ VPWR VPWR _379_/D _250_/D sky130_fd_sc_hd__fa_2
Xdadda_fa_4_98_0 dadda_fa_4_98_0/A dadda_fa_4_98_0/B dadda_fa_4_98_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_99_0/A dadda_fa_5_98_1/A sky130_fd_sc_hd__fa_1
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1305 U$$3972/A VGND VGND VPWR VPWR U$$3949/B sky130_fd_sc_hd__buf_6
Xfanout1316 U$$3835/A VGND VGND VPWR VPWR U$$3816/B sky130_fd_sc_hd__buf_6
Xfanout1327 input5/X VGND VGND VPWR VPWR U$$955/B sky130_fd_sc_hd__buf_8
XFILLER_78_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1338 input47/X VGND VGND VPWR VPWR U$$3474/B sky130_fd_sc_hd__clkbuf_4
Xfanout1349 input44/X VGND VGND VPWR VPWR U$$3425/A sky130_fd_sc_hd__buf_4
XFILLER_87_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout395 U$$904/A2 VGND VGND VPWR VPWR U$$876/A2 sky130_fd_sc_hd__buf_4
XU$$3107 U$$3107/A U$$3107/B VGND VGND VPWR VPWR U$$3107/X sky130_fd_sc_hd__xor2_1
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3118 U$$4486/B1 U$$3118/A2 U$$4353/A1 U$$3118/B2 VGND VGND VPWR VPWR U$$3119/A
+ sky130_fd_sc_hd__a22o_1
XU$$3129 U$$3129/A U$$3150/A VGND VGND VPWR VPWR U$$3129/X sky130_fd_sc_hd__xor2_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2406 U$$2406/A U$$2446/B VGND VGND VPWR VPWR U$$2406/X sky130_fd_sc_hd__xor2_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2417 U$$4196/B1 U$$2463/A2 U$$4198/B1 U$$2463/B2 VGND VGND VPWR VPWR U$$2418/A
+ sky130_fd_sc_hd__a22o_1
XU$$2428 U$$2428/A U$$2446/B VGND VGND VPWR VPWR U$$2428/X sky130_fd_sc_hd__xor2_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2439 U$$2576/A1 U$$2443/A2 U$$2576/B1 U$$2443/B2 VGND VGND VPWR VPWR U$$2440/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1705 U$$1705/A U$$1721/B VGND VGND VPWR VPWR U$$1705/X sky130_fd_sc_hd__xor2_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1716 U$$346/A1 U$$1720/A2 U$$2814/A1 U$$1720/B2 VGND VGND VPWR VPWR U$$1717/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1727 U$$1727/A U$$1727/B VGND VGND VPWR VPWR U$$1727/X sky130_fd_sc_hd__xor2_1
XFILLER_43_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1738 U$$3106/B1 U$$1774/A2 U$$3110/A1 U$$1774/B2 VGND VGND VPWR VPWR U$$1739/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1749 U$$1749/A U$$1761/B VGND VGND VPWR VPWR U$$1749/X sky130_fd_sc_hd__xor2_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_315_ _321_/CLK _315_/D VGND VGND VPWR VPWR _315_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_246_ _247_/CLK _246_/D VGND VGND VPWR VPWR _246_/Q sky130_fd_sc_hd__dfxtp_1
Xinput15 a[22] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput26 a[32] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_1
Xinput37 a[42] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
Xinput48 a[52] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput59 a[62] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_177_ _319_/CLK _177_/D VGND VGND VPWR VPWR _177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_62_5 dadda_fa_2_62_5/A dadda_fa_2_62_5/B dadda_fa_2_62_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_2/A dadda_fa_4_62_0/A sky130_fd_sc_hd__fa_2
XFILLER_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_55_4 dadda_fa_2_55_4/A dadda_fa_2_55_4/B dadda_fa_2_55_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_1/CIN dadda_fa_3_55_3/CIN sky130_fd_sc_hd__fa_1
XU$$4320 U$$4320/A U$$4322/B VGND VGND VPWR VPWR U$$4320/X sky130_fd_sc_hd__xor2_1
XU$$4331 U$$4331/A1 U$$4359/A2 U$$908/A1 U$$4359/B2 VGND VGND VPWR VPWR U$$4332/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3559_1821 VGND VGND VPWR VPWR U$$3559_1821/HI U$$3559/B1 sky130_fd_sc_hd__conb_1
XU$$4342 U$$4342/A U$$4350/B VGND VGND VPWR VPWR U$$4342/X sky130_fd_sc_hd__xor2_1
XU$$4353 U$$4353/A1 U$$4373/A2 U$$4353/B1 U$$4373/B2 VGND VGND VPWR VPWR U$$4354/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_48_3 dadda_fa_2_48_3/A dadda_fa_2_48_3/B dadda_fa_2_48_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_1/B dadda_fa_3_48_3/B sky130_fd_sc_hd__fa_1
XFILLER_38_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4364 U$$4364/A U$$4368/B VGND VGND VPWR VPWR U$$4364/X sky130_fd_sc_hd__xor2_1
XU$$3630 U$$4176/B1 U$$3640/A2 U$$3630/B1 U$$3640/B2 VGND VGND VPWR VPWR U$$3631/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4375 U$$4375/A1 U$$4381/A2 U$$4375/B1 U$$4381/B2 VGND VGND VPWR VPWR U$$4376/A
+ sky130_fd_sc_hd__a22o_1
XU$$4386 U$$4386/A VGND VGND VPWR VPWR U$$4386/Y sky130_fd_sc_hd__inv_1
XU$$3641 U$$3641/A U$$3641/B VGND VGND VPWR VPWR U$$3641/X sky130_fd_sc_hd__xor2_1
XFILLER_65_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4397 U$$4397/A U$$4397/B VGND VGND VPWR VPWR U$$4397/X sky130_fd_sc_hd__xor2_1
XFILLER_93_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3652 U$$4198/B1 U$$3682/A2 U$$4476/A1 U$$3682/B2 VGND VGND VPWR VPWR U$$3653/A
+ sky130_fd_sc_hd__a22o_1
XU$$3663 U$$3663/A U$$3681/B VGND VGND VPWR VPWR U$$3663/X sky130_fd_sc_hd__xor2_1
XU$$3674 U$$4359/A1 U$$3682/A2 U$$4359/B1 U$$3682/B2 VGND VGND VPWR VPWR U$$3675/A
+ sky130_fd_sc_hd__a22o_1
XU$$2940 U$$2940/A U$$3014/A VGND VGND VPWR VPWR U$$2940/X sky130_fd_sc_hd__xor2_1
XFILLER_52_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_18_1 dadda_fa_5_18_1/A dadda_fa_5_18_1/B dadda_fa_5_18_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_19_0/B dadda_fa_7_18_0/A sky130_fd_sc_hd__fa_1
XU$$3685 U$$3685/A U$$3695/B VGND VGND VPWR VPWR U$$3685/X sky130_fd_sc_hd__xor2_1
XU$$3696 U$$4107/A1 U$$3696/A2 U$$3696/B1 U$$3696/B2 VGND VGND VPWR VPWR U$$3697/A
+ sky130_fd_sc_hd__a22o_1
XU$$2951 U$$4456/B1 U$$3005/A2 U$$4049/A1 U$$3005/B2 VGND VGND VPWR VPWR U$$2952/A
+ sky130_fd_sc_hd__a22o_1
XU$$2962 U$$2962/A U$$2974/B VGND VGND VPWR VPWR U$$2962/X sky130_fd_sc_hd__xor2_1
XFILLER_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2973 U$$2973/A1 U$$2979/A2 U$$2973/B1 U$$2979/B2 VGND VGND VPWR VPWR U$$2974/A
+ sky130_fd_sc_hd__a22o_1
XU$$2984 U$$2984/A U$$2986/B VGND VGND VPWR VPWR U$$2984/X sky130_fd_sc_hd__xor2_1
XU$$2995 U$$3817/A1 U$$3005/A2 U$$3817/B1 U$$3005/B2 VGND VGND VPWR VPWR U$$2996/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_clk _201_/CLK VGND VGND VPWR VPWR _358_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$913 final_adder.U$$142/A final_adder.U$$851/X final_adder.U$$913/B1
+ VGND VGND VPWR VPWR final_adder.U$$913/X sky130_fd_sc_hd__a21o_1
XFILLER_84_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$935 final_adder.U$$164/A final_adder.U$$873/X final_adder.U$$935/B1
+ VGND VGND VPWR VPWR final_adder.U$$935/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_3 U$$1304/X U$$1437/X U$$1570/X VGND VGND VPWR VPWR dadda_fa_2_51_1/B
+ dadda_fa_2_50_4/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$957 final_adder.U$$186/A final_adder.U$$895/X final_adder.U$$957/B1
+ VGND VGND VPWR VPWR final_adder.U$$957/X sky130_fd_sc_hd__a21o_1
XU$$807 U$$944/A1 U$$807/A2 U$$944/B1 U$$807/B2 VGND VGND VPWR VPWR U$$808/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$979 final_adder.U$$208/A final_adder.U$$821/X final_adder.U$$979/B1
+ VGND VGND VPWR VPWR final_adder.U$$979/X sky130_fd_sc_hd__a21o_1
XU$$818 U$$818/A U$$820/B VGND VGND VPWR VPWR U$$818/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_43_2 U$$891/X U$$1024/X U$$1157/X VGND VGND VPWR VPWR dadda_fa_2_44_3/B
+ dadda_fa_2_43_5/B sky130_fd_sc_hd__fa_1
XU$$829 U$$829/A U$$875/B VGND VGND VPWR VPWR U$$829/X sky130_fd_sc_hd__xor2_1
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_20_1 dadda_fa_4_20_1/A dadda_fa_4_20_1/B dadda_fa_4_20_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_21_0/B dadda_fa_5_20_1/B sky130_fd_sc_hd__fa_1
XFILLER_25_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_13_0 U$$33/X U$$166/X U$$299/X VGND VGND VPWR VPWR dadda_fa_5_14_0/A dadda_fa_5_13_1/A
+ sky130_fd_sc_hd__fa_1
XFILLER_25_975 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1102 U$$54/A1 VGND VGND VPWR VPWR U$$465/A1 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_3_65_3 dadda_fa_3_65_3/A dadda_fa_3_65_3/B dadda_fa_3_65_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_1/B dadda_fa_4_65_2/CIN sky130_fd_sc_hd__fa_1
Xfanout1113 U$$874/A1 VGND VGND VPWR VPWR U$$50/B1 sky130_fd_sc_hd__buf_4
XFILLER_120_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1124 U$$3610/B1 VGND VGND VPWR VPWR U$$4434/A1 sky130_fd_sc_hd__buf_6
Xfanout1135 U$$4257/A1 VGND VGND VPWR VPWR U$$3296/B1 sky130_fd_sc_hd__buf_6
Xfanout1146 input75/X VGND VGND VPWR VPWR U$$4291/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_58_2 dadda_fa_3_58_2/A dadda_fa_3_58_2/B dadda_fa_3_58_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_1/A dadda_fa_4_58_2/B sky130_fd_sc_hd__fa_1
Xfanout1157 U$$4152/B1 VGND VGND VPWR VPWR U$$316/B1 sky130_fd_sc_hd__buf_4
Xfanout1168 U$$3189/B1 VGND VGND VPWR VPWR U$$997/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1179 U$$4422/A1 VGND VGND VPWR VPWR U$$3189/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_28_0 dadda_fa_6_28_0/A dadda_fa_6_28_0/B dadda_fa_6_28_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_29_0/B dadda_fa_7_28_0/CIN sky130_fd_sc_hd__fa_1
XU$$2203 U$$2203/A U$$2253/B VGND VGND VPWR VPWR U$$2203/X sky130_fd_sc_hd__xor2_1
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2214 U$$981/A1 U$$2272/A2 U$$981/B1 U$$2272/B2 VGND VGND VPWR VPWR U$$2215/A sky130_fd_sc_hd__a22o_1
XFILLER_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2225 U$$2225/A U$$2231/B VGND VGND VPWR VPWR U$$2225/X sky130_fd_sc_hd__xor2_1
XU$$2236 U$$2647/A1 U$$2252/A2 U$$46/A1 U$$2252/B2 VGND VGND VPWR VPWR U$$2237/A sky130_fd_sc_hd__a22o_1
XU$$1502 U$$4377/B1 U$$1502/A2 U$$4244/A1 U$$1502/B2 VGND VGND VPWR VPWR U$$1503/A
+ sky130_fd_sc_hd__a22o_1
XU$$2247 U$$2247/A U$$2249/B VGND VGND VPWR VPWR U$$2247/X sky130_fd_sc_hd__xor2_1
XFILLER_16_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2258 U$$66/A1 U$$2272/A2 U$$68/A1 U$$2272/B2 VGND VGND VPWR VPWR U$$2259/A sky130_fd_sc_hd__a22o_1
XU$$1513 U$$1513/A1 U$$1575/A2 U$$2748/A1 U$$1575/B2 VGND VGND VPWR VPWR U$$1514/A
+ sky130_fd_sc_hd__a22o_1
XU$$1524 U$$1524/A U$$1564/B VGND VGND VPWR VPWR U$$1524/X sky130_fd_sc_hd__xor2_1
XU$$2269 U$$2269/A U$$2269/B VGND VGND VPWR VPWR U$$2269/X sky130_fd_sc_hd__xor2_1
XFILLER_50_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1535 U$$576/A1 U$$1575/A2 U$$576/B1 U$$1575/B2 VGND VGND VPWR VPWR U$$1536/A sky130_fd_sc_hd__a22o_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1546 U$$1546/A U$$1584/B VGND VGND VPWR VPWR U$$1546/X sky130_fd_sc_hd__xor2_1
XU$$1557 U$$596/B1 U$$1563/A2 U$$598/B1 U$$1563/B2 VGND VGND VPWR VPWR U$$1558/A sky130_fd_sc_hd__a22o_1
XFILLER_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1568 U$$1568/A U$$1568/B VGND VGND VPWR VPWR U$$1568/X sky130_fd_sc_hd__xor2_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1579 U$$346/A1 U$$1621/A2 U$$2814/A1 U$$1621/B2 VGND VGND VPWR VPWR U$$1580/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2463_1803 VGND VGND VPWR VPWR U$$2463_1803/HI U$$2463/B1 sky130_fd_sc_hd__conb_1
XFILLER_30_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_229_ _358_/CLK _229_/D VGND VGND VPWR VPWR _229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_956 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_2 dadda_fa_2_60_2/A dadda_fa_2_60_2/B dadda_fa_2_60_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_1/A dadda_fa_3_60_3/A sky130_fd_sc_hd__fa_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$209 final_adder.U$$208/B final_adder.U$$979/B1 final_adder.U$$209/B1
+ VGND VGND VPWR VPWR final_adder.U$$209/X sky130_fd_sc_hd__a21o_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_53_1 dadda_fa_2_53_1/A dadda_fa_2_53_1/B dadda_fa_2_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_0/CIN dadda_fa_3_53_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1680 U$$2711/A1 VGND VGND VPWR VPWR fanout1680/X sky130_fd_sc_hd__buf_4
Xfanout1691 input11/X VGND VGND VPWR VPWR U$$1360/B sky130_fd_sc_hd__buf_6
Xdadda_fa_5_30_0 dadda_fa_5_30_0/A dadda_fa_5_30_0/B dadda_fa_5_30_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_31_0/A dadda_fa_6_30_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_46_0 U$$2759/X U$$2892/X U$$3025/X VGND VGND VPWR VPWR dadda_fa_3_47_0/B
+ dadda_fa_3_46_2/B sky130_fd_sc_hd__fa_1
XU$$4150 U$$4150/A1 U$$4240/A2 U$$4152/A1 U$$4240/B2 VGND VGND VPWR VPWR U$$4151/A
+ sky130_fd_sc_hd__a22o_1
XU$$4161 U$$4161/A U$$4175/B VGND VGND VPWR VPWR U$$4161/X sky130_fd_sc_hd__xor2_1
XU$$4172 U$$4307/B1 U$$4174/A2 U$$4174/A1 U$$4174/B2 VGND VGND VPWR VPWR U$$4173/A
+ sky130_fd_sc_hd__a22o_1
XU$$4183 U$$4183/A U$$4231/B VGND VGND VPWR VPWR U$$4183/X sky130_fd_sc_hd__xor2_1
XFILLER_92_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4194 U$$4331/A1 U$$4226/A2 U$$4196/A1 U$$4226/B2 VGND VGND VPWR VPWR U$$4195/A
+ sky130_fd_sc_hd__a22o_1
XU$$3460 U$$3460/A U$$3468/B VGND VGND VPWR VPWR U$$3460/X sky130_fd_sc_hd__xor2_1
XU$$3471 U$$4291/B1 U$$3471/A2 U$$4432/A1 U$$3471/B2 VGND VGND VPWR VPWR U$$3472/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3482 U$$3482/A U$$3482/B VGND VGND VPWR VPWR U$$3482/X sky130_fd_sc_hd__xor2_1
XU$$3493 U$$3628/B1 U$$3505/A2 U$$3630/B1 U$$3505/B2 VGND VGND VPWR VPWR U$$3494/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2770 U$$30/A1 U$$2856/A2 U$$32/A1 U$$2856/B2 VGND VGND VPWR VPWR U$$2771/A sky130_fd_sc_hd__a22o_1
XU$$2781 U$$2781/A U$$2811/B VGND VGND VPWR VPWR U$$2781/X sky130_fd_sc_hd__xor2_1
XU$$2792 U$$735/B1 U$$2798/A2 U$$602/A1 U$$2798/B2 VGND VGND VPWR VPWR U$$2793/A sky130_fd_sc_hd__a22o_1
XFILLER_21_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_75_2 dadda_fa_4_75_2/A dadda_fa_4_75_2/B dadda_fa_4_75_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_76_0/CIN dadda_fa_5_75_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_68_1 dadda_fa_4_68_1/A dadda_fa_4_68_1/B dadda_fa_4_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_69_0/B dadda_fa_5_68_1/B sky130_fd_sc_hd__fa_1
XFILLER_88_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput205 c[53] VGND VGND VPWR VPWR input205/X sky130_fd_sc_hd__buf_2
Xinput216 c[63] VGND VGND VPWR VPWR input216/X sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_7_45_0 dadda_fa_7_45_0/A dadda_fa_7_45_0/B dadda_fa_7_45_0/CIN VGND VGND
+ VPWR VPWR _342_/D _213_/D sky130_fd_sc_hd__fa_1
XFILLER_88_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput227 c[73] VGND VGND VPWR VPWR input227/X sky130_fd_sc_hd__buf_2
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput238 c[83] VGND VGND VPWR VPWR input238/X sky130_fd_sc_hd__dlymetal6s2s_1
Xdadda_ha_1_35_0 U$$77/X U$$210/X VGND VGND VPWR VPWR dadda_fa_2_36_5/B dadda_fa_3_35_0/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$710 final_adder.U$$710/A final_adder.U$$710/B VGND VGND VPWR VPWR
+ final_adder.U$$790/A sky130_fd_sc_hd__and2_1
Xinput249 c[93] VGND VGND VPWR VPWR input249/X sky130_fd_sc_hd__buf_2
Xfinal_adder.U$$721 final_adder.U$$720/B final_adder.U$$617/X final_adder.U$$601/X
+ VGND VGND VPWR VPWR final_adder.U$$721/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$743 final_adder.U$$742/B final_adder.U$$663/X final_adder.U$$631/X
+ VGND VGND VPWR VPWR final_adder.U$$743/X sky130_fd_sc_hd__a21o_1
XFILLER_57_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$754 final_adder.U$$786/B final_adder.U$$754/B VGND VGND VPWR VPWR
+ final_adder.U$$754/X sky130_fd_sc_hd__and2_1
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$765 final_adder.U$$764/B final_adder.U$$685/X final_adder.U$$653/X
+ VGND VGND VPWR VPWR final_adder.U$$765/X sky130_fd_sc_hd__a21o_1
XU$$604 U$$741/A1 U$$638/A2 U$$880/A1 U$$638/B2 VGND VGND VPWR VPWR U$$605/A sky130_fd_sc_hd__a22o_1
XFILLER_29_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$776 final_adder.U$$776/A final_adder.U$$776/B VGND VGND VPWR VPWR
+ final_adder.U$$776/X sky130_fd_sc_hd__and2_1
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$615 U$$615/A U$$639/B VGND VGND VPWR VPWR U$$615/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$787 final_adder.U$$786/B final_adder.U$$707/X final_adder.U$$675/X
+ VGND VGND VPWR VPWR final_adder.U$$787/X sky130_fd_sc_hd__a21o_1
XU$$626 U$$900/A1 U$$630/A2 U$$900/B1 U$$630/B2 VGND VGND VPWR VPWR U$$627/A sky130_fd_sc_hd__a22o_1
XFILLER_57_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$798 final_adder.U$$798/A final_adder.U$$798/B VGND VGND VPWR VPWR
+ final_adder.U$$798/X sky130_fd_sc_hd__and2_1
XU$$637 U$$637/A U$$637/B VGND VGND VPWR VPWR U$$637/X sky130_fd_sc_hd__xor2_1
XU$$648 U$$783/B1 U$$682/A2 U$$650/A1 U$$682/B2 VGND VGND VPWR VPWR U$$649/A sky130_fd_sc_hd__a22o_1
XU$$659 U$$659/A U$$669/B VGND VGND VPWR VPWR U$$659/X sky130_fd_sc_hd__xor2_1
XFILLER_16_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_916 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2189_1799 VGND VGND VPWR VPWR U$$2189_1799/HI U$$2189/B1 sky130_fd_sc_hd__conb_1
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_70_1 dadda_fa_3_70_1/A dadda_fa_3_70_1/B dadda_fa_3_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_0/CIN dadda_fa_4_70_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_63_0 dadda_fa_3_63_0/A dadda_fa_3_63_0/B dadda_fa_3_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_0/B dadda_fa_4_63_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2000 U$$3642/B1 U$$2046/A2 U$$3509/A1 U$$2046/B2 VGND VGND VPWR VPWR U$$2001/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2011 U$$2011/A U$$2053/B VGND VGND VPWR VPWR U$$2011/X sky130_fd_sc_hd__xor2_1
XU$$2022 U$$4486/B1 U$$2022/A2 U$$654/A1 U$$2022/B2 VGND VGND VPWR VPWR U$$2023/A
+ sky130_fd_sc_hd__a22o_1
XU$$2033 U$$2033/A U$$2043/B VGND VGND VPWR VPWR U$$2033/X sky130_fd_sc_hd__xor2_1
XFILLER_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2044 U$$2179/B1 U$$2044/A2 U$$2183/A1 U$$2044/B2 VGND VGND VPWR VPWR U$$2045/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2055 U$$2055/A VGND VGND VPWR VPWR U$$2055/Y sky130_fd_sc_hd__inv_1
XU$$1310 U$$1310/A U$$1320/B VGND VGND VPWR VPWR U$$1310/X sky130_fd_sc_hd__xor2_1
XU$$2066 U$$2066/A U$$2096/B VGND VGND VPWR VPWR U$$2066/X sky130_fd_sc_hd__xor2_1
XU$$1321 U$$773/A1 U$$1359/A2 U$$773/B1 U$$1359/B2 VGND VGND VPWR VPWR U$$1322/A sky130_fd_sc_hd__a22o_1
XU$$1332 U$$1332/A U$$1370/A VGND VGND VPWR VPWR U$$1332/X sky130_fd_sc_hd__xor2_1
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2077 U$$707/A1 U$$2107/A2 U$$709/A1 U$$2107/B2 VGND VGND VPWR VPWR U$$2078/A sky130_fd_sc_hd__a22o_1
XU$$2088 U$$2088/A U$$2096/B VGND VGND VPWR VPWR U$$2088/X sky130_fd_sc_hd__xor2_1
XU$$1343 U$$521/A1 U$$1359/A2 U$$521/B1 U$$1359/B2 VGND VGND VPWR VPWR U$$1344/A sky130_fd_sc_hd__a22o_1
XU$$1354 U$$1354/A U$$1358/B VGND VGND VPWR VPWR U$$1354/X sky130_fd_sc_hd__xor2_1
XU$$2099 U$$866/A1 U$$2107/A2 U$$868/A1 U$$2107/B2 VGND VGND VPWR VPWR U$$2100/A sky130_fd_sc_hd__a22o_1
XU$$1365 U$$406/A1 U$$1367/A2 U$$406/B1 U$$1367/B2 VGND VGND VPWR VPWR U$$1366/A sky130_fd_sc_hd__a22o_1
XU$$1376 U$$1376/A1 U$$1452/A2 U$$828/B1 U$$1452/B2 VGND VGND VPWR VPWR U$$1377/A
+ sky130_fd_sc_hd__a22o_1
XU$$1387 U$$1387/A U$$1433/B VGND VGND VPWR VPWR U$$1387/X sky130_fd_sc_hd__xor2_1
XFILLER_149_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1398 U$$850/A1 U$$1426/A2 U$$989/A1 U$$1426/B2 VGND VGND VPWR VPWR U$$1399/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_7_120_0 dadda_fa_7_120_0/A dadda_fa_7_120_0/B dadda_fa_7_120_0/CIN VGND
+ VGND VPWR VPWR _417_/D _288_/D sky130_fd_sc_hd__fa_1
XFILLER_148_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_85_1 dadda_fa_5_85_1/A dadda_fa_5_85_1/B dadda_fa_5_85_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_86_0/B dadda_fa_7_85_0/A sky130_fd_sc_hd__fa_2
XFILLER_7_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_78_0 dadda_fa_5_78_0/A dadda_fa_5_78_0/B dadda_fa_5_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_79_0/A dadda_fa_6_78_0/CIN sky130_fd_sc_hd__fa_1
Xfanout906 U$$1202/B2 VGND VGND VPWR VPWR U$$1230/B2 sky130_fd_sc_hd__buf_6
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout917 U$$74/B2 VGND VGND VPWR VPWR U$$80/B2 sky130_fd_sc_hd__buf_2
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_77_8 input231/X dadda_fa_1_77_8/B dadda_fa_1_77_8/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_78_3/A dadda_fa_3_77_0/A sky130_fd_sc_hd__fa_1
Xfanout928 U$$4389/X VGND VGND VPWR VPWR U$$4502/B2 sky130_fd_sc_hd__clkbuf_2
Xfanout939 U$$2480/A1 VGND VGND VPWR VPWR U$$2754/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$50 _346_/Q _218_/Q VGND VGND VPWR VPWR final_adder.U$$975/B1 final_adder.U$$204/A
+ sky130_fd_sc_hd__ha_2
XFILLER_81_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$61 _357_/Q _229_/Q VGND VGND VPWR VPWR final_adder.U$$195/B1 final_adder.U$$194/B
+ sky130_fd_sc_hd__ha_1
XFILLER_54_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3290 U$$3425/A VGND VGND VPWR VPWR U$$3290/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$72 _368_/Q _240_/Q VGND VGND VPWR VPWR final_adder.U$$953/B1 final_adder.U$$182/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$83 _379_/Q _251_/Q VGND VGND VPWR VPWR final_adder.U$$173/B1 final_adder.U$$172/B
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$94 _390_/Q _262_/Q VGND VGND VPWR VPWR final_adder.U$$931/B1 final_adder.U$$160/A
+ sky130_fd_sc_hd__ha_1
XFILLER_16_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_80_0 dadda_fa_4_80_0/A dadda_fa_4_80_0/B dadda_fa_4_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_81_0/A dadda_fa_5_80_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_101_3 dadda_fa_3_101_3/A dadda_fa_3_101_3/B dadda_fa_3_101_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_102_1/B dadda_fa_4_101_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$540 final_adder.U$$548/B final_adder.U$$540/B VGND VGND VPWR VPWR
+ final_adder.U$$660/B sky130_fd_sc_hd__and2_1
XFILLER_29_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$551 final_adder.U$$550/B final_adder.U$$435/X final_adder.U$$427/X
+ VGND VGND VPWR VPWR final_adder.U$$551/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$562 final_adder.U$$570/B final_adder.U$$562/B VGND VGND VPWR VPWR
+ final_adder.U$$682/B sky130_fd_sc_hd__and2_1
XU$$401 U$$401/A U$$411/A VGND VGND VPWR VPWR U$$401/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_108_0 dadda_fa_6_108_0/A dadda_fa_6_108_0/B dadda_fa_6_108_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_109_0/B dadda_fa_7_108_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$573 final_adder.U$$572/B final_adder.U$$457/X final_adder.U$$449/X
+ VGND VGND VPWR VPWR final_adder.U$$573/X sky130_fd_sc_hd__a21o_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$412 U$$412/A VGND VGND VPWR VPWR U$$414/B sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$584 final_adder.U$$592/B final_adder.U$$584/B VGND VGND VPWR VPWR
+ final_adder.U$$704/B sky130_fd_sc_hd__and2_1
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$423 U$$12/A1 U$$447/A2 U$$14/A1 U$$447/B2 VGND VGND VPWR VPWR U$$424/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$595 final_adder.U$$594/B final_adder.U$$479/X final_adder.U$$471/X
+ VGND VGND VPWR VPWR final_adder.U$$595/X sky130_fd_sc_hd__a21o_1
XFILLER_72_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$434 U$$434/A U$$448/B VGND VGND VPWR VPWR U$$434/X sky130_fd_sc_hd__xor2_1
XU$$445 U$$32/B1 U$$447/A2 U$$447/A1 U$$447/B2 VGND VGND VPWR VPWR U$$446/A sky130_fd_sc_hd__a22o_1
XU$$456 U$$456/A U$$498/B VGND VGND VPWR VPWR U$$456/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_28_3 dadda_fa_3_28_3/A dadda_fa_3_28_3/B dadda_fa_3_28_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_29_1/B dadda_fa_4_28_2/CIN sky130_fd_sc_hd__fa_1
XU$$467 U$$56/A1 U$$501/A2 U$$56/B1 U$$501/B2 VGND VGND VPWR VPWR U$$468/A sky130_fd_sc_hd__a22o_1
XU$$478 U$$478/A U$$480/B VGND VGND VPWR VPWR U$$478/X sky130_fd_sc_hd__xor2_1
XU$$489 U$$900/A1 U$$497/A2 U$$900/B1 U$$497/B2 VGND VGND VPWR VPWR U$$490/A sky130_fd_sc_hd__a22o_1
XFILLER_32_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_95_0 dadda_fa_6_95_0/A dadda_fa_6_95_0/B dadda_fa_6_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_96_0/B dadda_fa_7_95_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_30_3 U$$1264/X U$$1397/X U$$1530/X VGND VGND VPWR VPWR dadda_fa_3_31_2/A
+ dadda_fa_3_30_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_91_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$990 U$$990/A U$$990/B VGND VGND VPWR VPWR U$$990/X sky130_fd_sc_hd__xor2_1
XFILLER_51_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1140 U$$44/A1 U$$1174/A2 U$$46/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1141/A sky130_fd_sc_hd__a22o_1
XU$$1151 U$$1151/A U$$1195/B VGND VGND VPWR VPWR U$$1151/X sky130_fd_sc_hd__xor2_1
XU$$1162 U$$64/B1 U$$1194/A2 U$$66/B1 U$$1194/B2 VGND VGND VPWR VPWR U$$1163/A sky130_fd_sc_hd__a22o_1
XFILLER_50_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1173 U$$1173/A U$$1175/B VGND VGND VPWR VPWR U$$1173/X sky130_fd_sc_hd__xor2_1
XU$$1184 U$$773/A1 U$$1226/A2 U$$773/B1 U$$1226/B2 VGND VGND VPWR VPWR U$$1185/A sky130_fd_sc_hd__a22o_1
XU$$1195 U$$1195/A U$$1195/B VGND VGND VPWR VPWR U$$1195/X sky130_fd_sc_hd__xor2_1
XFILLER_137_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_82_6 U$$3629/X U$$3762/X U$$3895/X VGND VGND VPWR VPWR dadda_fa_2_83_3/B
+ dadda_fa_2_82_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_49_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout703 U$$4115/X VGND VGND VPWR VPWR U$$4244/B2 sky130_fd_sc_hd__buf_6
Xfanout714 U$$3978/X VGND VGND VPWR VPWR U$$4107/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_160_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout725 U$$3924/B2 VGND VGND VPWR VPWR U$$3966/B2 sky130_fd_sc_hd__buf_2
Xdadda_fa_1_75_5 U$$3615/X U$$3748/X U$$3881/X VGND VGND VPWR VPWR dadda_fa_2_76_2/A
+ dadda_fa_2_75_5/A sky130_fd_sc_hd__fa_1
Xfanout736 U$$3644/B2 VGND VGND VPWR VPWR U$$3640/B2 sky130_fd_sc_hd__buf_4
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout747 U$$3439/B2 VGND VGND VPWR VPWR U$$3523/B2 sky130_fd_sc_hd__buf_6
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout758 U$$3422/B2 VGND VGND VPWR VPWR U$$3418/B2 sky130_fd_sc_hd__buf_2
Xfanout769 U$$3156/X VGND VGND VPWR VPWR U$$3257/B2 sky130_fd_sc_hd__clkbuf_8
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_4 U$$4133/X U$$4266/X U$$4399/X VGND VGND VPWR VPWR dadda_fa_2_69_1/CIN
+ dadda_fa_2_68_4/CIN sky130_fd_sc_hd__fa_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_38_2 dadda_fa_4_38_2/A dadda_fa_4_38_2/B dadda_fa_4_38_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_39_0/CIN dadda_fa_5_38_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3696_1823 VGND VGND VPWR VPWR U$$3696_1823/HI U$$3696/B1 sky130_fd_sc_hd__conb_1
Xdadda_fa_0_63_3 U$$1330/X U$$1463/X U$$1596/X VGND VGND VPWR VPWR dadda_fa_1_64_6/B
+ dadda_fa_1_63_8/B sky130_fd_sc_hd__fa_1
XFILLER_76_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_40_2 dadda_fa_3_40_2/A dadda_fa_3_40_2/B dadda_fa_3_40_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_1/A dadda_fa_4_40_2/B sky130_fd_sc_hd__fa_1
XFILLER_58_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$370 final_adder.U$$372/B final_adder.U$$370/B VGND VGND VPWR VPWR
+ final_adder.U$$496/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$381 final_adder.U$$378/A final_adder.U$$255/X final_adder.U$$253/X
+ VGND VGND VPWR VPWR final_adder.U$$381/X sky130_fd_sc_hd__a21o_2
XU$$220 U$$220/A U$$220/B VGND VGND VPWR VPWR U$$220/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_33_1 dadda_fa_3_33_1/A dadda_fa_3_33_1/B dadda_fa_3_33_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_34_0/CIN dadda_fa_4_33_2/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$392 final_adder.U$$396/B final_adder.U$$392/B VGND VGND VPWR VPWR
+ final_adder.U$$516/B sky130_fd_sc_hd__and2_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$231 U$$94/A1 U$$271/A2 U$$96/A1 U$$271/B2 VGND VGND VPWR VPWR U$$232/A sky130_fd_sc_hd__a22o_1
XFILLER_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$242 U$$242/A U$$254/B VGND VGND VPWR VPWR U$$242/X sky130_fd_sc_hd__xor2_1
XFILLER_55_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_10_0 dadda_fa_6_10_0/A dadda_fa_6_10_0/B dadda_fa_6_10_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_11_0/B dadda_fa_7_10_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_26_0 U$$1123/X U$$1256/X U$$1389/X VGND VGND VPWR VPWR dadda_fa_4_27_0/B
+ dadda_fa_4_26_1/CIN sky130_fd_sc_hd__fa_1
XU$$253 U$$253/A1 U$$253/A2 U$$253/B1 U$$253/B2 VGND VGND VPWR VPWR U$$254/A sky130_fd_sc_hd__a22o_1
XU$$264 U$$264/A U$$274/A VGND VGND VPWR VPWR U$$264/X sky130_fd_sc_hd__xor2_1
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$275 U$$275/A VGND VGND VPWR VPWR U$$277/B sky130_fd_sc_hd__inv_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$286 U$$12/A1 U$$312/A2 U$$14/A1 U$$312/B2 VGND VGND VPWR VPWR U$$287/A sky130_fd_sc_hd__a22o_1
XFILLER_60_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$297 U$$297/A U$$313/B VGND VGND VPWR VPWR U$$297/X sky130_fd_sc_hd__xor2_1
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3 U$$3/A U$$3/B VGND VGND VPWR VPWR U$$3/X sky130_fd_sc_hd__and2_1
XFILLER_127_931 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput306 output306/A VGND VGND VPWR VPWR o[29] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_5 dadda_fa_2_92_5/A dadda_fa_2_92_5/B dadda_fa_2_92_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_93_2/A dadda_fa_4_92_0/A sky130_fd_sc_hd__fa_1
XFILLER_154_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput317 output317/A VGND VGND VPWR VPWR o[39] sky130_fd_sc_hd__buf_2
Xoutput328 output328/A VGND VGND VPWR VPWR o[49] sky130_fd_sc_hd__buf_2
Xoutput339 output339/A VGND VGND VPWR VPWR o[59] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_85_4 dadda_fa_2_85_4/A dadda_fa_2_85_4/B dadda_fa_2_85_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_1/CIN dadda_fa_3_85_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_78_3 dadda_fa_2_78_3/A dadda_fa_2_78_3/B dadda_fa_2_78_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_1/B dadda_fa_3_78_3/B sky130_fd_sc_hd__fa_1
XFILLER_45_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1040 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_48_1 dadda_fa_5_48_1/A dadda_fa_5_48_1/B dadda_fa_5_48_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_49_0/B dadda_fa_7_48_0/A sky130_fd_sc_hd__fa_1
XFILLER_67_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_101_2 U$$3401/X U$$3534/X U$$3667/X VGND VGND VPWR VPWR dadda_fa_3_102_2/B
+ dadda_fa_3_101_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_32_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_122_1 input154/X dadda_fa_5_122_1/B dadda_ha_4_122_0/SUM VGND VGND VPWR
+ VPWR dadda_fa_6_123_0/B dadda_fa_7_122_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_115_0 dadda_fa_5_115_0/A dadda_fa_5_115_0/B dadda_fa_5_115_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_116_0/A dadda_fa_6_115_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_80_3 U$$2295/X U$$2428/X U$$2561/X VGND VGND VPWR VPWR dadda_fa_2_81_1/CIN
+ dadda_fa_2_80_4/B sky130_fd_sc_hd__fa_1
Xfanout500 U$$3306/A2 VGND VGND VPWR VPWR U$$3422/A2 sky130_fd_sc_hd__buf_4
Xfanout511 U$$3072/A2 VGND VGND VPWR VPWR U$$3066/A2 sky130_fd_sc_hd__buf_4
Xfanout1509 input128/X VGND VGND VPWR VPWR U$$985/A1 sky130_fd_sc_hd__buf_6
XFILLER_120_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout522 U$$2977/A2 VGND VGND VPWR VPWR U$$2979/A2 sky130_fd_sc_hd__buf_4
Xfanout533 U$$346/A2 VGND VGND VPWR VPWR U$$340/A2 sky130_fd_sc_hd__buf_2
Xdadda_fa_1_73_2 U$$2680/X U$$2813/X U$$2946/X VGND VGND VPWR VPWR dadda_fa_2_74_1/A
+ dadda_fa_2_73_4/A sky130_fd_sc_hd__fa_1
Xfanout544 U$$2744/X VGND VGND VPWR VPWR U$$2812/A2 sky130_fd_sc_hd__buf_4
Xfanout555 fanout561/X VGND VGND VPWR VPWR U$$2574/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_4_50_1 dadda_fa_4_50_1/A dadda_fa_4_50_1/B dadda_fa_4_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_51_0/B dadda_fa_5_50_1/B sky130_fd_sc_hd__fa_1
XFILLER_59_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_66_1 U$$2932/X U$$3065/X U$$3198/X VGND VGND VPWR VPWR dadda_fa_2_67_0/CIN
+ dadda_fa_2_66_3/CIN sky130_fd_sc_hd__fa_1
Xfanout566 U$$2463/A2 VGND VGND VPWR VPWR U$$2415/A2 sky130_fd_sc_hd__clkbuf_8
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout577 U$$2196/X VGND VGND VPWR VPWR U$$2320/A2 sky130_fd_sc_hd__buf_4
XFILLER_101_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_2_100_4 U$$4064/X U$$4197/X VGND VGND VPWR VPWR dadda_fa_3_101_2/CIN dadda_fa_4_100_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout588 U$$2014/A2 VGND VGND VPWR VPWR U$$1980/A2 sky130_fd_sc_hd__clkbuf_4
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_43_0 dadda_fa_4_43_0/A dadda_fa_4_43_0/B dadda_fa_4_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_44_0/A dadda_fa_5_43_1/A sky130_fd_sc_hd__fa_1
Xfanout599 U$$1915/A2 VGND VGND VPWR VPWR U$$1909/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_59_0 U$$1588/X U$$1721/X U$$1854/X VGND VGND VPWR VPWR dadda_fa_2_60_0/B
+ dadda_fa_2_59_3/B sky130_fd_sc_hd__fa_1
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_400_ _402_/CLK _400_/D VGND VGND VPWR VPWR _400_/Q sky130_fd_sc_hd__dfxtp_1
XU$$1909 U$$2183/A1 U$$1909/A2 U$$4512/B1 U$$1909/B2 VGND VGND VPWR VPWR U$$1910/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_331_ _344_/CLK _331_/D VGND VGND VPWR VPWR _331_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_262_ _408_/CLK _262_/D VGND VGND VPWR VPWR _262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_193_ _321_/CLK _193_/D VGND VGND VPWR VPWR _193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_931 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_95_3 dadda_fa_3_95_3/A dadda_fa_3_95_3/B dadda_fa_3_95_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_1/B dadda_fa_4_95_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_6_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_88_2 dadda_fa_3_88_2/A dadda_fa_3_88_2/B dadda_fa_3_88_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_1/A dadda_fa_4_88_2/B sky130_fd_sc_hd__fa_1
Xdadda_ha_0_55_1 U$$516/X U$$649/X VGND VGND VPWR VPWR dadda_fa_1_56_8/A dadda_fa_2_55_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_58_0 dadda_fa_6_58_0/A dadda_fa_6_58_0/B dadda_fa_6_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_59_0/B dadda_fa_7_58_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_110_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4502 U$$4502/A1 U$$4388/X U$$4504/A1 U$$4502/B2 VGND VGND VPWR VPWR U$$4503/A
+ sky130_fd_sc_hd__a22o_1
XU$$4513 U$$4513/A U$$4513/B VGND VGND VPWR VPWR U$$4513/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_61_0 U$$129/X U$$262/X U$$395/X VGND VGND VPWR VPWR dadda_fa_1_62_5/CIN
+ dadda_fa_1_61_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_65_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3801 U$$4484/B1 U$$3833/A2 U$$4488/A1 U$$3833/B2 VGND VGND VPWR VPWR U$$3802/A
+ sky130_fd_sc_hd__a22o_1
XU$$16 U$$16/A1 U$$8/A2 U$$18/A1 U$$8/B2 VGND VGND VPWR VPWR U$$17/A sky130_fd_sc_hd__a22o_1
XU$$3812 U$$3812/A U$$3816/B VGND VGND VPWR VPWR U$$3812/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_117_2 U$$4497/X input148/X dadda_fa_4_117_2/CIN VGND VGND VPWR VPWR dadda_fa_5_118_0/CIN
+ dadda_fa_5_117_1/CIN sky130_fd_sc_hd__fa_1
XU$$3823 U$$3960/A1 U$$3833/A2 U$$4508/B1 U$$3833/B2 VGND VGND VPWR VPWR U$$3824/A
+ sky130_fd_sc_hd__a22o_1
XU$$27 U$$27/A U$$49/B VGND VGND VPWR VPWR U$$27/X sky130_fd_sc_hd__xor2_1
XFILLER_64_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$38 U$$38/A1 U$$74/A2 U$$40/A1 U$$74/B2 VGND VGND VPWR VPWR U$$39/A sky130_fd_sc_hd__a22o_1
XU$$3834 U$$3834/A U$$3835/A VGND VGND VPWR VPWR U$$3834/X sky130_fd_sc_hd__xor2_1
XU$$49 U$$49/A U$$49/B VGND VGND VPWR VPWR U$$49/X sky130_fd_sc_hd__xor2_1
XFILLER_80_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3845 U$$3845/A U$$3925/B VGND VGND VPWR VPWR U$$3845/X sky130_fd_sc_hd__xor2_1
XU$$3856 U$$4265/B1 U$$3892/A2 U$$4132/A1 U$$3892/B2 VGND VGND VPWR VPWR U$$3857/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3867 U$$3867/A U$$3867/B VGND VGND VPWR VPWR U$$3867/X sky130_fd_sc_hd__xor2_1
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3878 U$$4152/A1 U$$3924/A2 U$$4152/B1 U$$3924/B2 VGND VGND VPWR VPWR U$$3879/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3889 U$$3889/A U$$3907/B VGND VGND VPWR VPWR U$$3889/X sky130_fd_sc_hd__xor2_1
XFILLER_61_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_976 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_90_2 U$$4044/X U$$4177/X U$$4310/X VGND VGND VPWR VPWR dadda_fa_3_91_1/A
+ dadda_fa_3_90_3/A sky130_fd_sc_hd__fa_1
XFILLER_115_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_83_1 input238/X dadda_fa_2_83_1/B dadda_fa_2_83_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_84_0/CIN dadda_fa_3_83_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_60_0 dadda_fa_5_60_0/A dadda_fa_5_60_0/B dadda_fa_5_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_61_0/A dadda_fa_6_60_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_76_0 dadda_fa_2_76_0/A dadda_fa_2_76_0/B dadda_fa_2_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_0/B dadda_fa_3_76_2/B sky130_fd_sc_hd__fa_1
XFILLER_28_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_52_7 U$$3170/X U$$3303/X U$$3436/X VGND VGND VPWR VPWR dadda_fa_2_53_2/CIN
+ dadda_fa_2_52_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_78_0_1942 VGND VGND VPWR VPWR dadda_ha_0_78_0/A dadda_ha_0_78_0_1942/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_98_1 dadda_fa_4_98_1/A dadda_fa_4_98_1/B dadda_fa_4_98_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_99_0/B dadda_fa_5_98_1/B sky130_fd_sc_hd__fa_1
XFILLER_152_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_75_0 dadda_fa_7_75_0/A dadda_fa_7_75_0/B dadda_fa_7_75_0/CIN VGND VGND
+ VPWR VPWR _372_/D _243_/D sky130_fd_sc_hd__fa_1
XFILLER_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1306 U$$3972/A VGND VGND VPWR VPWR U$$3961/B sky130_fd_sc_hd__clkbuf_4
Xfanout1317 U$$3792/B VGND VGND VPWR VPWR U$$3835/A sky130_fd_sc_hd__buf_6
Xfanout1328 U$$3607/B VGND VGND VPWR VPWR U$$3601/B sky130_fd_sc_hd__buf_6
Xfanout1339 U$$3562/A VGND VGND VPWR VPWR U$$3506/B sky130_fd_sc_hd__buf_6
XFILLER_87_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout385 U$$999/A2 VGND VGND VPWR VPWR U$$997/A2 sky130_fd_sc_hd__buf_4
XFILLER_74_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout396 U$$904/A2 VGND VGND VPWR VPWR U$$910/A2 sky130_fd_sc_hd__buf_2
XU$$3108 U$$3243/B1 U$$3108/A2 U$$3110/A1 U$$3108/B2 VGND VGND VPWR VPWR U$$3109/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3119 U$$3119/A U$$3119/B VGND VGND VPWR VPWR U$$3119/X sky130_fd_sc_hd__xor2_1
XFILLER_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2407 U$$3775/B1 U$$2407/A2 U$$902/A1 U$$2407/B2 VGND VGND VPWR VPWR U$$2408/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2418 U$$2418/A U$$2456/B VGND VGND VPWR VPWR U$$2418/X sky130_fd_sc_hd__xor2_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2429 U$$2840/A1 U$$2443/A2 U$$2840/B1 U$$2443/B2 VGND VGND VPWR VPWR U$$2430/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1706 U$$882/B1 U$$1720/A2 U$$747/B1 U$$1720/B2 VGND VGND VPWR VPWR U$$1707/A sky130_fd_sc_hd__a22o_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1717 U$$1717/A U$$1721/B VGND VGND VPWR VPWR U$$1717/X sky130_fd_sc_hd__xor2_1
XU$$1728 U$$3370/B1 U$$1774/A2 U$$632/B1 U$$1774/B2 VGND VGND VPWR VPWR U$$1729/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1739 U$$1739/A U$$1741/B VGND VGND VPWR VPWR U$$1739/X sky130_fd_sc_hd__xor2_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_314_ _321_/CLK _314_/D VGND VGND VPWR VPWR _314_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_245_ _375_/CLK _245_/D VGND VGND VPWR VPWR _245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput16 a[23] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__clkbuf_4
Xinput27 a[33] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_1
Xinput38 a[43] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_4
X_176_ _321_/CLK _176_/D VGND VGND VPWR VPWR _176_/Q sky130_fd_sc_hd__dfxtp_1
Xinput49 a[53] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_93_0 dadda_fa_3_93_0/A dadda_fa_3_93_0/B dadda_fa_3_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_0/B dadda_fa_4_93_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4310 U$$4310/A U$$4383/A VGND VGND VPWR VPWR U$$4310/X sky130_fd_sc_hd__xor2_1
XFILLER_93_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4321 U$$4456/B1 U$$4325/A2 U$$4460/A1 U$$4325/B2 VGND VGND VPWR VPWR U$$4322/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_55_5 dadda_fa_2_55_5/A dadda_fa_2_55_5/B dadda_fa_2_55_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_2/A dadda_fa_4_55_0/A sky130_fd_sc_hd__fa_1
XFILLER_42_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4332 U$$4332/A U$$4360/B VGND VGND VPWR VPWR U$$4332/X sky130_fd_sc_hd__xor2_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4343 U$$4478/B1 U$$4349/A2 U$$4345/A1 U$$4349/B2 VGND VGND VPWR VPWR U$$4344/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4354 U$$4354/A U$$4368/B VGND VGND VPWR VPWR U$$4354/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_48_4 dadda_fa_2_48_4/A dadda_fa_2_48_4/B dadda_fa_2_48_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_1/CIN dadda_fa_3_48_3/CIN sky130_fd_sc_hd__fa_1
XU$$3620 U$$4440/B1 U$$3644/A2 U$$4307/A1 U$$3644/B2 VGND VGND VPWR VPWR U$$3621/A
+ sky130_fd_sc_hd__a22o_1
XU$$4365 U$$4365/A1 U$$4373/A2 U$$4365/B1 U$$4373/B2 VGND VGND VPWR VPWR U$$4366/A
+ sky130_fd_sc_hd__a22o_1
XU$$3631 U$$3631/A U$$3641/B VGND VGND VPWR VPWR U$$3631/X sky130_fd_sc_hd__xor2_1
XU$$4376 U$$4376/A U$$4383/A VGND VGND VPWR VPWR U$$4376/X sky130_fd_sc_hd__xor2_1
XU$$4387 U$$4387/A U$$4387/B VGND VGND VPWR VPWR U$$4387/X sky130_fd_sc_hd__and2_1
XU$$3642 U$$3642/A1 U$$3644/A2 U$$3642/B1 U$$3644/B2 VGND VGND VPWR VPWR U$$3643/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4398 U$$4398/A1 U$$4388/X U$$4400/A1 U$$4428/B2 VGND VGND VPWR VPWR U$$4399/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3653 U$$3653/A U$$3681/B VGND VGND VPWR VPWR U$$3653/X sky130_fd_sc_hd__xor2_1
XU$$3664 U$$4484/B1 U$$3692/A2 U$$4349/B1 U$$3692/B2 VGND VGND VPWR VPWR U$$3665/A
+ sky130_fd_sc_hd__a22o_1
XU$$2930 U$$2930/A U$$2974/B VGND VGND VPWR VPWR U$$2930/X sky130_fd_sc_hd__xor2_1
XU$$3675 U$$3675/A U$$3698/A VGND VGND VPWR VPWR U$$3675/X sky130_fd_sc_hd__xor2_1
XU$$2941 U$$612/A1 U$$2991/A2 U$$612/B1 U$$2991/B2 VGND VGND VPWR VPWR U$$2942/A sky130_fd_sc_hd__a22o_1
XU$$3686 U$$4234/A1 U$$3692/A2 U$$4234/B1 U$$3692/B2 VGND VGND VPWR VPWR U$$3687/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3697 U$$3697/A U$$3698/A VGND VGND VPWR VPWR U$$3697/X sky130_fd_sc_hd__xor2_1
XU$$2952 U$$2952/A U$$3004/B VGND VGND VPWR VPWR U$$2952/X sky130_fd_sc_hd__xor2_1
XU$$2963 U$$3372/B1 U$$2979/A2 U$$3239/A1 U$$2979/B2 VGND VGND VPWR VPWR U$$2964/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2974 U$$2974/A U$$2974/B VGND VGND VPWR VPWR U$$2974/X sky130_fd_sc_hd__xor2_1
XU$$2985 U$$4353/B1 U$$3011/A2 U$$4220/A1 U$$3011/B2 VGND VGND VPWR VPWR U$$2986/A
+ sky130_fd_sc_hd__a22o_1
XU$$2996 U$$2996/A U$$3004/B VGND VGND VPWR VPWR U$$2996/X sky130_fd_sc_hd__xor2_1
XFILLER_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_1_44_5 U$$2090/X U$$2223/X VGND VGND VPWR VPWR dadda_fa_2_45_4/A dadda_fa_3_44_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_102_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$903 final_adder.U$$132/A final_adder.U$$841/X final_adder.U$$903/B1
+ VGND VGND VPWR VPWR final_adder.U$$903/X sky130_fd_sc_hd__a21o_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$925 final_adder.U$$154/A final_adder.U$$863/X final_adder.U$$925/B1
+ VGND VGND VPWR VPWR final_adder.U$$925/X sky130_fd_sc_hd__a21o_1
XFILLER_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$947 final_adder.U$$176/A final_adder.U$$885/X final_adder.U$$947/B1
+ VGND VGND VPWR VPWR final_adder.U$$947/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_4 U$$1703/X U$$1836/X U$$1969/X VGND VGND VPWR VPWR dadda_fa_2_51_1/CIN
+ dadda_fa_2_50_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$808 U$$808/A U$$822/A VGND VGND VPWR VPWR U$$808/X sky130_fd_sc_hd__xor2_1
XFILLER_83_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$969 final_adder.U$$198/A final_adder.U$$811/X final_adder.U$$969/B1
+ VGND VGND VPWR VPWR final_adder.U$$969/X sky130_fd_sc_hd__a21o_1
XFILLER_56_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$819 U$$956/A1 U$$819/A2 U$$819/B1 U$$819/B2 VGND VGND VPWR VPWR U$$820/A sky130_fd_sc_hd__a22o_1
XFILLER_113_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_43_3 U$$1290/X U$$1423/X U$$1556/X VGND VGND VPWR VPWR dadda_fa_2_44_3/CIN
+ dadda_fa_2_43_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_37_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_20_2 dadda_fa_4_20_2/A dadda_fa_4_20_2/B dadda_ha_3_20_3/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_21_0/CIN dadda_fa_5_20_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_71_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_13_1 U$$432/X U$$565/X U$$698/X VGND VGND VPWR VPWR dadda_fa_5_14_0/B
+ dadda_fa_5_13_1/B sky130_fd_sc_hd__fa_1
XFILLER_25_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_889 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1103 U$$602/A1 VGND VGND VPWR VPWR U$$54/A1 sky130_fd_sc_hd__buf_4
XFILLER_154_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1114 input79/X VGND VGND VPWR VPWR U$$874/A1 sky130_fd_sc_hd__buf_6
Xfanout1125 input78/X VGND VGND VPWR VPWR U$$3610/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1136 input76/X VGND VGND VPWR VPWR U$$4257/A1 sky130_fd_sc_hd__buf_4
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1147 U$$183/A1 VGND VGND VPWR VPWR U$$46/A1 sky130_fd_sc_hd__buf_4
Xfanout1158 input74/X VGND VGND VPWR VPWR U$$4152/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_58_3 dadda_fa_3_58_3/A dadda_fa_3_58_3/B dadda_fa_3_58_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_1/B dadda_fa_4_58_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1169 U$$3189/B1 VGND VGND VPWR VPWR U$$999/A1 sky130_fd_sc_hd__buf_4
XFILLER_102_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2204 U$$697/A1 U$$2248/A2 U$$697/B1 U$$2248/B2 VGND VGND VPWR VPWR U$$2205/A sky130_fd_sc_hd__a22o_1
XU$$2215 U$$2215/A U$$2231/B VGND VGND VPWR VPWR U$$2215/X sky130_fd_sc_hd__xor2_1
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2226 U$$856/A1 U$$2254/A2 U$$3322/B1 U$$2254/B2 VGND VGND VPWR VPWR U$$2227/A
+ sky130_fd_sc_hd__a22o_1
XU$$2237 U$$2237/A U$$2249/B VGND VGND VPWR VPWR U$$2237/X sky130_fd_sc_hd__xor2_1
XU$$1503 U$$1503/A U$$1507/A VGND VGND VPWR VPWR U$$1503/X sky130_fd_sc_hd__xor2_1
XU$$2248 U$$878/A1 U$$2248/A2 U$$878/B1 U$$2248/B2 VGND VGND VPWR VPWR U$$2249/A sky130_fd_sc_hd__a22o_1
XU$$2259 U$$2259/A U$$2269/B VGND VGND VPWR VPWR U$$2259/X sky130_fd_sc_hd__xor2_1
XU$$1514 U$$1514/A U$$1570/B VGND VGND VPWR VPWR U$$1514/X sky130_fd_sc_hd__xor2_1
XU$$1525 U$$2758/A1 U$$1563/A2 U$$2758/B1 U$$1563/B2 VGND VGND VPWR VPWR U$$1526/A
+ sky130_fd_sc_hd__a22o_1
XU$$1536 U$$1536/A U$$1570/B VGND VGND VPWR VPWR U$$1536/X sky130_fd_sc_hd__xor2_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1547 U$$40/A1 U$$1575/A2 U$$40/B1 U$$1575/B2 VGND VGND VPWR VPWR U$$1548/A sky130_fd_sc_hd__a22o_1
XU$$1558 U$$1558/A U$$1564/B VGND VGND VPWR VPWR U$$1558/X sky130_fd_sc_hd__xor2_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1569 U$$882/B1 U$$1587/A2 U$$747/B1 U$$1587/B2 VGND VGND VPWR VPWR U$$1570/A sky130_fd_sc_hd__a22o_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_228_ _358_/CLK _228_/D VGND VGND VPWR VPWR _228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_3 dadda_fa_2_60_3/A dadda_fa_2_60_3/B dadda_fa_2_60_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_1/B dadda_fa_3_60_3/B sky130_fd_sc_hd__fa_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_53_2 dadda_fa_2_53_2/A dadda_fa_2_53_2/B dadda_fa_2_53_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_1/A dadda_fa_3_53_3/A sky130_fd_sc_hd__fa_1
XFILLER_111_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1670 U$$4494/A1 VGND VGND VPWR VPWR U$$4492/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1681 input110/X VGND VGND VPWR VPWR U$$2711/A1 sky130_fd_sc_hd__buf_4
Xfanout1692 U$$3030/A1 VGND VGND VPWR VPWR U$$2891/B1 sky130_fd_sc_hd__clkbuf_4
XU$$4140 U$$4414/A1 U$$4190/A2 U$$4416/A1 U$$4190/B2 VGND VGND VPWR VPWR U$$4141/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_30_1 dadda_fa_5_30_1/A dadda_fa_5_30_1/B dadda_fa_5_30_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_31_0/B dadda_fa_7_30_0/A sky130_fd_sc_hd__fa_1
XU$$4151 U$$4151/A U$$4231/B VGND VGND VPWR VPWR U$$4151/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_46_1 U$$3158/X U$$3196/B input197/X VGND VGND VPWR VPWR dadda_fa_3_47_0/CIN
+ dadda_fa_3_46_2/CIN sky130_fd_sc_hd__fa_1
XU$$4162 U$$4162/A1 U$$4174/A2 U$$4162/B1 U$$4174/B2 VGND VGND VPWR VPWR U$$4163/A
+ sky130_fd_sc_hd__a22o_1
XU$$4173 U$$4173/A U$$4175/B VGND VGND VPWR VPWR U$$4173/X sky130_fd_sc_hd__xor2_1
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_23_0 dadda_fa_5_23_0/A dadda_fa_5_23_0/B dadda_fa_5_23_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_24_0/A dadda_fa_6_23_0/CIN sky130_fd_sc_hd__fa_2
XU$$4184 U$$4456/B1 U$$4224/A2 U$$4460/A1 U$$4224/B2 VGND VGND VPWR VPWR U$$4185/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3450 U$$3450/A U$$3468/B VGND VGND VPWR VPWR U$$3450/X sky130_fd_sc_hd__xor2_1
XU$$4195 U$$4195/A U$$4215/B VGND VGND VPWR VPWR U$$4195/X sky130_fd_sc_hd__xor2_1
XU$$3461 U$$3870/B1 U$$3471/A2 U$$4420/B1 U$$3471/B2 VGND VGND VPWR VPWR U$$3462/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_39_0 U$$1149/X U$$1282/X U$$1415/X VGND VGND VPWR VPWR dadda_fa_3_40_0/B
+ dadda_fa_3_39_2/B sky130_fd_sc_hd__fa_1
XFILLER_53_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3472 U$$3472/A U$$3474/B VGND VGND VPWR VPWR U$$3472/X sky130_fd_sc_hd__xor2_1
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3483 U$$3618/B1 U$$3557/A2 U$$4444/A1 U$$3557/B2 VGND VGND VPWR VPWR U$$3484/A
+ sky130_fd_sc_hd__a22o_1
XU$$3494 U$$3494/A U$$3506/B VGND VGND VPWR VPWR U$$3494/X sky130_fd_sc_hd__xor2_1
XU$$2760 U$$2897/A1 U$$2798/A2 U$$2897/B1 U$$2798/B2 VGND VGND VPWR VPWR U$$2761/A
+ sky130_fd_sc_hd__a22o_1
XU$$2771 U$$2771/A U$$2811/B VGND VGND VPWR VPWR U$$2771/X sky130_fd_sc_hd__xor2_1
XU$$2782 U$$40/B1 U$$2856/A2 U$$316/B1 U$$2856/B2 VGND VGND VPWR VPWR U$$2783/A sky130_fd_sc_hd__a22o_1
XFILLER_80_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2793 U$$2793/A U$$2799/B VGND VGND VPWR VPWR U$$2793/X sky130_fd_sc_hd__xor2_1
XFILLER_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_68_2 dadda_fa_4_68_2/A dadda_fa_4_68_2/B dadda_fa_4_68_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_69_0/CIN dadda_fa_5_68_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput206 c[54] VGND VGND VPWR VPWR input206/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput217 c[64] VGND VGND VPWR VPWR input217/X sky130_fd_sc_hd__clkbuf_1
Xinput228 c[74] VGND VGND VPWR VPWR input228/X sky130_fd_sc_hd__buf_2
Xinput239 c[84] VGND VGND VPWR VPWR input239/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$700 final_adder.U$$716/B final_adder.U$$700/B VGND VGND VPWR VPWR
+ final_adder.U$$780/A sky130_fd_sc_hd__and2_1
XFILLER_69_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$711 final_adder.U$$710/B final_adder.U$$607/X final_adder.U$$591/X
+ VGND VGND VPWR VPWR final_adder.U$$711/X sky130_fd_sc_hd__a21o_1
XFILLER_124_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_38_0 dadda_fa_7_38_0/A dadda_fa_7_38_0/B dadda_fa_7_38_0/CIN VGND VGND
+ VPWR VPWR _335_/D _206_/D sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$733 final_adder.U$$716/A final_adder.U$$505/X final_adder.U$$613/X
+ VGND VGND VPWR VPWR final_adder.U$$733/X sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$744 final_adder.U$$776/B final_adder.U$$744/B VGND VGND VPWR VPWR
+ final_adder.U$$744/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$755 final_adder.U$$754/B final_adder.U$$675/X final_adder.U$$643/X
+ VGND VGND VPWR VPWR final_adder.U$$755/X sky130_fd_sc_hd__a21o_1
XFILLER_57_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$766 final_adder.U$$798/B final_adder.U$$766/B VGND VGND VPWR VPWR
+ final_adder.U$$766/X sky130_fd_sc_hd__and2_1
XFILLER_17_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$605 U$$605/A U$$639/B VGND VGND VPWR VPWR U$$605/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$777 final_adder.U$$776/B final_adder.U$$697/X final_adder.U$$665/X
+ VGND VGND VPWR VPWR final_adder.U$$777/X sky130_fd_sc_hd__a21o_1
XU$$616 U$$616/A1 U$$636/A2 U$$892/A1 U$$636/B2 VGND VGND VPWR VPWR U$$617/A sky130_fd_sc_hd__a22o_1
XFILLER_72_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$788 final_adder.U$$788/A final_adder.U$$788/B VGND VGND VPWR VPWR
+ final_adder.U$$788/X sky130_fd_sc_hd__and2_1
XU$$627 U$$627/A U$$631/B VGND VGND VPWR VPWR U$$627/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_41_0 U$$89/X U$$222/X U$$355/X VGND VGND VPWR VPWR dadda_fa_2_42_3/B dadda_fa_2_41_5/A
+ sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$799 final_adder.U$$798/B final_adder.U$$719/X final_adder.U$$687/X
+ VGND VGND VPWR VPWR final_adder.U$$799/X sky130_fd_sc_hd__a21o_1
XU$$638 U$$773/B1 U$$638/A2 U$$640/A1 U$$638/B2 VGND VGND VPWR VPWR U$$639/A sky130_fd_sc_hd__a22o_1
XU$$649 U$$649/A U$$684/A VGND VGND VPWR VPWR U$$649/X sky130_fd_sc_hd__xor2_1
XFILLER_140_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_928 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_70_2 dadda_fa_3_70_2/A dadda_fa_3_70_2/B dadda_fa_3_70_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_1/A dadda_fa_4_70_2/B sky130_fd_sc_hd__fa_1
XFILLER_3_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$5_1907 VGND VGND VPWR VPWR U$$5_1907/HI U$$5/A2 sky130_fd_sc_hd__conb_1
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_63_1 dadda_fa_3_63_1/A dadda_fa_3_63_1/B dadda_fa_3_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_0/CIN dadda_fa_4_63_2/A sky130_fd_sc_hd__fa_1
XFILLER_79_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_40_0 dadda_fa_6_40_0/A dadda_fa_6_40_0/B dadda_fa_6_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_41_0/B dadda_fa_7_40_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_56_0 dadda_fa_3_56_0/A dadda_fa_3_56_0/B dadda_fa_3_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_0/B dadda_fa_4_56_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2001 U$$2001/A U$$2031/B VGND VGND VPWR VPWR U$$2001/X sky130_fd_sc_hd__xor2_1
XU$$2012 U$$916/A1 U$$2014/A2 U$$918/A1 U$$2014/B2 VGND VGND VPWR VPWR U$$2013/A sky130_fd_sc_hd__a22o_1
XFILLER_35_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2023 U$$2023/A U$$2053/B VGND VGND VPWR VPWR U$$2023/X sky130_fd_sc_hd__xor2_1
XU$$2034 U$$2443/B1 U$$2044/A2 U$$2310/A1 U$$2044/B2 VGND VGND VPWR VPWR U$$2035/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1300 U$$1300/A U$$1300/B VGND VGND VPWR VPWR U$$1300/X sky130_fd_sc_hd__xor2_1
XU$$2045 U$$2045/A U$$2055/A VGND VGND VPWR VPWR U$$2045/X sky130_fd_sc_hd__xor2_1
XFILLER_62_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2056 input24/X VGND VGND VPWR VPWR U$$2058/B sky130_fd_sc_hd__inv_1
XFILLER_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1311 U$$78/A1 U$$1311/A2 U$$80/A1 U$$1311/B2 VGND VGND VPWR VPWR U$$1312/A sky130_fd_sc_hd__a22o_1
XU$$1322 U$$1322/A U$$1360/B VGND VGND VPWR VPWR U$$1322/X sky130_fd_sc_hd__xor2_1
XU$$2067 U$$3298/B1 U$$2107/A2 U$$2480/A1 U$$2107/B2 VGND VGND VPWR VPWR U$$2068/A
+ sky130_fd_sc_hd__a22o_1
XU$$1333 U$$2840/A1 U$$1367/A2 U$$2840/B1 U$$1367/B2 VGND VGND VPWR VPWR U$$1334/A
+ sky130_fd_sc_hd__a22o_1
XU$$2078 U$$2078/A U$$2106/B VGND VGND VPWR VPWR U$$2078/X sky130_fd_sc_hd__xor2_1
XU$$2089 U$$993/A1 U$$2097/A2 U$$995/A1 U$$2097/B2 VGND VGND VPWR VPWR U$$2090/A sky130_fd_sc_hd__a22o_1
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1344 U$$1344/A U$$1358/B VGND VGND VPWR VPWR U$$1344/X sky130_fd_sc_hd__xor2_1
XU$$1355 U$$120/B1 U$$1359/A2 U$$946/A1 U$$1359/B2 VGND VGND VPWR VPWR U$$1356/A sky130_fd_sc_hd__a22o_1
XU$$1366 U$$1366/A U$$1370/A VGND VGND VPWR VPWR U$$1366/X sky130_fd_sc_hd__xor2_1
XU$$1377 U$$1377/A U$$1415/B VGND VGND VPWR VPWR U$$1377/X sky130_fd_sc_hd__xor2_1
XFILLER_31_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1388 U$$2758/A1 U$$1426/A2 U$$2758/B1 U$$1426/B2 VGND VGND VPWR VPWR U$$1389/A
+ sky130_fd_sc_hd__a22o_1
XU$$1399 U$$1399/A U$$1427/B VGND VGND VPWR VPWR U$$1399/X sky130_fd_sc_hd__xor2_1
XFILLER_90_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_113_0 dadda_fa_7_113_0/A dadda_fa_7_113_0/B dadda_fa_7_113_0/CIN VGND
+ VGND VPWR VPWR _410_/D _281_/D sky130_fd_sc_hd__fa_1
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_78_1 dadda_fa_5_78_1/A dadda_fa_5_78_1/B dadda_fa_5_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_79_0/B dadda_fa_7_78_0/A sky130_fd_sc_hd__fa_2
XFILLER_135_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout907 U$$1170/B2 VGND VGND VPWR VPWR U$$1174/B2 sky130_fd_sc_hd__buf_4
Xfanout918 U$$120/B2 VGND VGND VPWR VPWR U$$74/B2 sky130_fd_sc_hd__clkbuf_4
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 fanout938/X VGND VGND VPWR VPWR U$$499/A1 sky130_fd_sc_hd__buf_4
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$40 _336_/Q _208_/Q VGND VGND VPWR VPWR final_adder.U$$985/B1 final_adder.U$$214/A
+ sky130_fd_sc_hd__ha_1
XFILLER_26_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$51 _347_/Q _219_/Q VGND VGND VPWR VPWR final_adder.U$$205/B1 final_adder.U$$204/B
+ sky130_fd_sc_hd__ha_2
XU$$3280 U$$3280/A U$$3284/B VGND VGND VPWR VPWR U$$3280/X sky130_fd_sc_hd__xor2_1
XU$$3291 U$$3425/A U$$3291/B VGND VGND VPWR VPWR U$$3291/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$62 _358_/Q _230_/Q VGND VGND VPWR VPWR final_adder.U$$963/B1 final_adder.U$$192/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$73 _369_/Q _241_/Q VGND VGND VPWR VPWR final_adder.U$$183/B1 final_adder.U$$182/B
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$84 _380_/Q _252_/Q VGND VGND VPWR VPWR final_adder.U$$941/B1 final_adder.U$$170/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$95 _391_/Q _263_/Q VGND VGND VPWR VPWR final_adder.U$$161/B1 final_adder.U$$160/B
+ sky130_fd_sc_hd__ha_1
XU$$2590 U$$946/A1 U$$2598/A2 U$$948/A1 U$$2598/B2 VGND VGND VPWR VPWR U$$2591/A sky130_fd_sc_hd__a22o_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_80_1 dadda_fa_4_80_1/A dadda_fa_4_80_1/B dadda_fa_4_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_81_0/B dadda_fa_5_80_1/B sky130_fd_sc_hd__fa_1
XFILLER_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_73_0 dadda_fa_4_73_0/A dadda_fa_4_73_0/B dadda_fa_4_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_74_0/A dadda_fa_5_73_1/A sky130_fd_sc_hd__fa_1
XFILLER_116_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_89_0 U$$1780/Y U$$1914/X U$$2047/X VGND VGND VPWR VPWR dadda_fa_2_90_3/CIN
+ dadda_fa_2_89_5/A sky130_fd_sc_hd__fa_1
XFILLER_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$530 final_adder.U$$538/B final_adder.U$$530/B VGND VGND VPWR VPWR
+ final_adder.U$$650/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$541 final_adder.U$$540/B final_adder.U$$425/X final_adder.U$$417/X
+ VGND VGND VPWR VPWR final_adder.U$$541/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$552 final_adder.U$$560/B final_adder.U$$552/B VGND VGND VPWR VPWR
+ final_adder.U$$672/B sky130_fd_sc_hd__and2_1
XFILLER_29_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$563 final_adder.U$$562/B final_adder.U$$447/X final_adder.U$$439/X
+ VGND VGND VPWR VPWR final_adder.U$$563/X sky130_fd_sc_hd__a21o_1
XU$$402 U$$539/A1 U$$406/A2 U$$539/B1 U$$406/B2 VGND VGND VPWR VPWR U$$403/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$574 final_adder.U$$582/B final_adder.U$$574/B VGND VGND VPWR VPWR
+ final_adder.U$$694/B sky130_fd_sc_hd__and2_1
XU$$413 U$$536/B VGND VGND VPWR VPWR U$$413/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$585 final_adder.U$$584/B final_adder.U$$469/X final_adder.U$$461/X
+ VGND VGND VPWR VPWR final_adder.U$$585/X sky130_fd_sc_hd__a21o_1
XU$$424 U$$424/A U$$448/B VGND VGND VPWR VPWR U$$424/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$596 final_adder.U$$604/B final_adder.U$$596/B VGND VGND VPWR VPWR
+ final_adder.U$$716/B sky130_fd_sc_hd__and2_1
XU$$435 U$$709/A1 U$$505/A2 U$$709/B1 U$$505/B2 VGND VGND VPWR VPWR U$$436/A sky130_fd_sc_hd__a22o_1
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$446 U$$446/A U$$448/B VGND VGND VPWR VPWR U$$446/X sky130_fd_sc_hd__xor2_1
XU$$457 U$$729/B1 U$$497/A2 U$$596/A1 U$$497/B2 VGND VGND VPWR VPWR U$$458/A sky130_fd_sc_hd__a22o_1
XU$$468 U$$468/A U$$504/B VGND VGND VPWR VPWR U$$468/X sky130_fd_sc_hd__xor2_1
XU$$479 U$$479/A1 U$$479/A2 U$$479/B1 U$$479/B2 VGND VGND VPWR VPWR U$$480/A sky130_fd_sc_hd__a22o_1
XFILLER_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2052_1797 VGND VGND VPWR VPWR U$$2052_1797/HI U$$2052/B1 sky130_fd_sc_hd__conb_1
XFILLER_157_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_88_0 dadda_fa_6_88_0/A dadda_fa_6_88_0/B dadda_fa_6_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_89_0/B dadda_fa_7_88_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_126_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_78_0 dadda_ha_0_78_0/A U$$1094/X VGND VGND VPWR VPWR dadda_fa_2_79_0/A
+ dadda_fa_2_78_0/A sky130_fd_sc_hd__ha_1
XFILLER_158_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$980 U$$980/A U$$980/B VGND VGND VPWR VPWR U$$980/X sky130_fd_sc_hd__xor2_1
XU$$991 U$$991/A1 U$$997/A2 U$$993/A1 U$$997/B2 VGND VGND VPWR VPWR U$$992/A sky130_fd_sc_hd__a22o_1
XU$$1130 U$$993/A1 U$$1164/A2 U$$995/A1 U$$1164/B2 VGND VGND VPWR VPWR U$$1131/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_92_0_1929 VGND VGND VPWR VPWR dadda_fa_1_92_0/A dadda_fa_1_92_0_1929/LO
+ sky130_fd_sc_hd__conb_1
XU$$1141 U$$1141/A U$$1175/B VGND VGND VPWR VPWR U$$1141/X sky130_fd_sc_hd__xor2_1
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1152 U$$465/B1 U$$1194/A2 U$$58/A1 U$$1194/B2 VGND VGND VPWR VPWR U$$1153/A sky130_fd_sc_hd__a22o_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1163 U$$1163/A U$$1163/B VGND VGND VPWR VPWR U$$1163/X sky130_fd_sc_hd__xor2_1
XFILLER_50_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1174 U$$78/A1 U$$1174/A2 U$$80/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1175/A sky130_fd_sc_hd__a22o_1
XU$$1185 U$$1185/A U$$1227/B VGND VGND VPWR VPWR U$$1185/X sky130_fd_sc_hd__xor2_1
XU$$1196 U$$2840/A1 U$$1230/A2 U$$2840/B1 U$$1230/B2 VGND VGND VPWR VPWR U$$1197/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_90_0 dadda_fa_5_90_0/A dadda_fa_5_90_0/B dadda_fa_5_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_91_0/A dadda_fa_6_90_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout704 U$$4190/B2 VGND VGND VPWR VPWR U$$4240/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout715 U$$4057/B2 VGND VGND VPWR VPWR U$$4081/B2 sky130_fd_sc_hd__buf_4
Xfanout726 U$$3841/X VGND VGND VPWR VPWR U$$3924/B2 sky130_fd_sc_hd__buf_6
Xfanout737 U$$3567/X VGND VGND VPWR VPWR U$$3644/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_75_6 U$$4014/X U$$4147/X U$$4280/X VGND VGND VPWR VPWR dadda_fa_2_76_2/B
+ dadda_fa_2_75_5/B sky130_fd_sc_hd__fa_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 U$$3439/B2 VGND VGND VPWR VPWR U$$3549/B2 sky130_fd_sc_hd__buf_4
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout759 U$$3306/B2 VGND VGND VPWR VPWR U$$3422/B2 sky130_fd_sc_hd__buf_4
XFILLER_140_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_5 input221/X dadda_fa_1_68_5/B dadda_fa_1_68_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_69_2/A dadda_fa_2_68_5/A sky130_fd_sc_hd__fa_1
XFILLER_58_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_120_0 dadda_fa_6_120_0/A dadda_fa_6_120_0/B dadda_fa_6_120_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_121_0/B dadda_fa_7_120_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_63_4 U$$1729/X U$$1862/X U$$1995/X VGND VGND VPWR VPWR dadda_fa_1_64_6/CIN
+ dadda_fa_1_63_8/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_40_3 dadda_fa_3_40_3/A dadda_fa_3_40_3/B dadda_fa_3_40_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_1/B dadda_fa_4_40_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_92_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$360 final_adder.U$$362/B final_adder.U$$360/B VGND VGND VPWR VPWR
+ final_adder.U$$486/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$371 final_adder.U$$370/B final_adder.U$$245/X final_adder.U$$243/X
+ VGND VGND VPWR VPWR final_adder.U$$371/X sky130_fd_sc_hd__a21o_1
XU$$210 U$$210/A U$$210/B VGND VGND VPWR VPWR U$$210/X sky130_fd_sc_hd__xor2_1
XU$$221 U$$84/A1 U$$229/A2 U$$86/A1 U$$229/B2 VGND VGND VPWR VPWR U$$222/A sky130_fd_sc_hd__a22o_1
XFILLER_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_33_2 dadda_fa_3_33_2/A dadda_fa_3_33_2/B dadda_fa_3_33_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_34_1/A dadda_fa_4_33_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$393 final_adder.U$$392/B final_adder.U$$271/X final_adder.U$$267/X
+ VGND VGND VPWR VPWR final_adder.U$$393/X sky130_fd_sc_hd__a21o_1
XU$$232 U$$232/A U$$273/A VGND VGND VPWR VPWR U$$232/X sky130_fd_sc_hd__xor2_1
XFILLER_44_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$243 U$$654/A1 U$$253/A2 U$$654/B1 U$$253/B2 VGND VGND VPWR VPWR U$$244/A sky130_fd_sc_hd__a22o_1
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$254 U$$254/A U$$254/B VGND VGND VPWR VPWR U$$254/X sky130_fd_sc_hd__xor2_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_26_1 U$$1522/X U$$1655/X U$$1788/X VGND VGND VPWR VPWR dadda_fa_4_27_0/CIN
+ dadda_fa_4_26_2/A sky130_fd_sc_hd__fa_1
XU$$265 U$$539/A1 U$$271/A2 U$$539/B1 U$$271/B2 VGND VGND VPWR VPWR U$$266/A sky130_fd_sc_hd__a22o_1
XFILLER_55_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$276 U$$411/A VGND VGND VPWR VPWR U$$276/Y sky130_fd_sc_hd__inv_1
XFILLER_55_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$287 U$$287/A U$$313/B VGND VGND VPWR VPWR U$$287/X sky130_fd_sc_hd__xor2_1
XFILLER_72_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$298 U$$24/A1 U$$312/A2 U$$26/A1 U$$312/B2 VGND VGND VPWR VPWR U$$299/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_19_0 U$$45/X U$$178/X U$$311/X VGND VGND VPWR VPWR dadda_fa_4_20_0/CIN
+ dadda_fa_4_19_2/A sky130_fd_sc_hd__fa_1
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4 U$$2/Y U$$1/A U$$4/A3 U$$3/X U$$0/Y VGND VGND VPWR VPWR U$$4/X sky130_fd_sc_hd__a32o_1
XFILLER_127_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput307 output307/A VGND VGND VPWR VPWR o[2] sky130_fd_sc_hd__buf_2
XFILLER_160_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput318 output318/A VGND VGND VPWR VPWR o[3] sky130_fd_sc_hd__buf_2
Xoutput329 output329/A VGND VGND VPWR VPWR o[4] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_85_5 dadda_fa_2_85_5/A dadda_fa_2_85_5/B dadda_fa_2_85_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_2/A dadda_fa_4_85_0/A sky130_fd_sc_hd__fa_2
XFILLER_113_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_78_4 dadda_fa_2_78_4/A dadda_fa_2_78_4/B dadda_fa_2_78_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_1/CIN dadda_fa_3_78_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_45_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_101_3 U$$3800/X U$$3933/X U$$4066/X VGND VGND VPWR VPWR dadda_fa_3_102_2/CIN
+ dadda_fa_4_101_0/A sky130_fd_sc_hd__fa_1
XFILLER_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_115_1 dadda_fa_5_115_1/A dadda_fa_5_115_1/B dadda_fa_5_115_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_116_0/B dadda_fa_7_115_0/A sky130_fd_sc_hd__fa_1
XFILLER_118_954 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_108_0 dadda_fa_5_108_0/A dadda_fa_5_108_0/B dadda_fa_5_108_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_109_0/A dadda_fa_6_108_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_80_4 U$$2694/X U$$2827/X U$$2960/X VGND VGND VPWR VPWR dadda_fa_2_81_2/A
+ dadda_fa_2_80_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout501 U$$3292/X VGND VGND VPWR VPWR U$$3306/A2 sky130_fd_sc_hd__buf_4
Xfanout512 U$$3112/A2 VGND VGND VPWR VPWR U$$3072/A2 sky130_fd_sc_hd__buf_4
Xfanout523 U$$2881/X VGND VGND VPWR VPWR U$$2977/A2 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_1_73_3 U$$3079/X U$$3212/X U$$3345/X VGND VGND VPWR VPWR dadda_fa_2_74_1/B
+ dadda_fa_2_73_4/B sky130_fd_sc_hd__fa_1
XFILLER_76_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout534 U$$338/A2 VGND VGND VPWR VPWR U$$346/A2 sky130_fd_sc_hd__clkbuf_2
Xfanout545 U$$2667/A2 VGND VGND VPWR VPWR U$$2665/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_4_50_2 dadda_fa_4_50_2/A dadda_fa_4_50_2/B dadda_fa_4_50_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_51_0/CIN dadda_fa_5_50_1/CIN sky130_fd_sc_hd__fa_1
Xfanout556 fanout561/X VGND VGND VPWR VPWR U$$2578/A2 sky130_fd_sc_hd__buf_2
Xdadda_fa_1_66_2 U$$3331/X U$$3464/X U$$3597/X VGND VGND VPWR VPWR dadda_fa_2_67_1/A
+ dadda_fa_2_66_4/A sky130_fd_sc_hd__fa_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout567 U$$2463/A2 VGND VGND VPWR VPWR U$$2413/A2 sky130_fd_sc_hd__buf_4
Xfanout578 U$$2139/A2 VGND VGND VPWR VPWR U$$2097/A2 sky130_fd_sc_hd__buf_4
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout589 U$$2022/A2 VGND VGND VPWR VPWR U$$2014/A2 sky130_fd_sc_hd__buf_4
XFILLER_101_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_43_1 dadda_fa_4_43_1/A dadda_fa_4_43_1/B dadda_fa_4_43_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_44_0/B dadda_fa_5_43_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_59_1 U$$1987/X U$$2120/X U$$2253/X VGND VGND VPWR VPWR dadda_fa_2_60_0/CIN
+ dadda_fa_2_59_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_7_20_0 dadda_fa_7_20_0/A dadda_fa_7_20_0/B dadda_fa_7_20_0/CIN VGND VGND
+ VPWR VPWR _317_/D _188_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_36_0 dadda_fa_4_36_0/A dadda_fa_4_36_0/B dadda_fa_4_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_37_0/A dadda_fa_5_36_1/A sky130_fd_sc_hd__fa_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_330_ _344_/CLK _330_/D VGND VGND VPWR VPWR _330_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_261_ _391_/CLK _261_/D VGND VGND VPWR VPWR _261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_192_ _328_/CLK _192_/D VGND VGND VPWR VPWR _192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_88_3 dadda_fa_3_88_3/A dadda_fa_3_88_3/B dadda_fa_3_88_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_1/B dadda_fa_4_88_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_2_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4431_1863 VGND VGND VPWR VPWR U$$4431_1863/HI U$$4431/B sky130_fd_sc_hd__conb_1
XFILLER_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4503 U$$4503/A U$$4503/B VGND VGND VPWR VPWR U$$4503/X sky130_fd_sc_hd__xor2_1
XU$$4514 U$$4514/A1 U$$4388/X U$$4516/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4515/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_0_61_1 U$$528/X U$$661/X U$$794/X VGND VGND VPWR VPWR dadda_fa_1_62_6/A
+ dadda_fa_1_61_8/A sky130_fd_sc_hd__fa_1
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3802 U$$3802/A U$$3816/B VGND VGND VPWR VPWR U$$3802/X sky130_fd_sc_hd__xor2_1
XU$$17 U$$17/A U$$9/B VGND VGND VPWR VPWR U$$17/X sky130_fd_sc_hd__xor2_1
XU$$3813 U$$3948/B1 U$$3825/A2 U$$3815/A1 U$$3825/B2 VGND VGND VPWR VPWR U$$3814/A
+ sky130_fd_sc_hd__a22o_1
XU$$28 U$$28/A1 U$$80/A2 U$$30/A1 U$$80/B2 VGND VGND VPWR VPWR U$$29/A sky130_fd_sc_hd__a22o_1
XFILLER_18_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3824 U$$3824/A U$$3828/B VGND VGND VPWR VPWR U$$3824/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_54_0 U$$115/X U$$248/X U$$381/X VGND VGND VPWR VPWR dadda_fa_1_55_8/A
+ dadda_fa_1_54_8/CIN sky130_fd_sc_hd__fa_1
XU$$39 U$$39/A U$$77/B VGND VGND VPWR VPWR U$$39/X sky130_fd_sc_hd__xor2_1
XU$$3835 U$$3835/A VGND VGND VPWR VPWR U$$3835/Y sky130_fd_sc_hd__inv_1
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3846 U$$3846/A1 U$$3872/A2 U$$3846/B1 U$$3872/B2 VGND VGND VPWR VPWR U$$3847/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4507_1901 VGND VGND VPWR VPWR U$$4507_1901/HI U$$4507/B sky130_fd_sc_hd__conb_1
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$190 final_adder.U$$190/A final_adder.U$$190/B VGND VGND VPWR VPWR
+ final_adder.U$$318/B sky130_fd_sc_hd__and2_1
XU$$3857 U$$3857/A U$$3867/B VGND VGND VPWR VPWR U$$3857/X sky130_fd_sc_hd__xor2_1
XU$$3868 U$$854/A1 U$$3872/A2 U$$3870/A1 U$$3872/B2 VGND VGND VPWR VPWR U$$3869/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3879 U$$3879/A U$$3925/B VGND VGND VPWR VPWR U$$3879/X sky130_fd_sc_hd__xor2_1
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_90_3 U$$4443/X input246/X dadda_fa_2_90_3/CIN VGND VGND VPWR VPWR dadda_fa_3_91_1/B
+ dadda_fa_3_90_3/B sky130_fd_sc_hd__fa_1
XFILLER_126_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_83_2 dadda_fa_2_83_2/A dadda_fa_2_83_2/B dadda_fa_2_83_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_1/A dadda_fa_3_83_3/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_60_1 dadda_fa_5_60_1/A dadda_fa_5_60_1/B dadda_fa_5_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_61_0/B dadda_fa_7_60_0/A sky130_fd_sc_hd__fa_2
XFILLER_87_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_76_1 dadda_fa_2_76_1/A dadda_fa_2_76_1/B dadda_fa_2_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_0/CIN dadda_fa_3_76_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_53_0 dadda_fa_5_53_0/A dadda_fa_5_53_0/B dadda_fa_5_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_54_0/A dadda_fa_6_53_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_69_0 dadda_fa_2_69_0/A dadda_fa_2_69_0/B dadda_fa_2_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_0/B dadda_fa_3_69_2/B sky130_fd_sc_hd__fa_1
XFILLER_110_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_52_8 U$$3569/X U$$3615/B input204/X VGND VGND VPWR VPWR dadda_fa_2_53_3/A
+ dadda_fa_3_52_0/A sky130_fd_sc_hd__fa_2
XU$$134_1785 VGND VGND VPWR VPWR U$$134_1785/HI U$$134/B1 sky130_fd_sc_hd__conb_1
XFILLER_52_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_98_2 dadda_fa_4_98_2/A dadda_fa_4_98_2/B dadda_fa_4_98_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_99_0/CIN dadda_fa_5_98_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_139_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_68_0 dadda_fa_7_68_0/A dadda_fa_7_68_0/B dadda_fa_7_68_0/CIN VGND VGND
+ VPWR VPWR _365_/D _236_/D sky130_fd_sc_hd__fa_1
XFILLER_160_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1307 fanout1309/X VGND VGND VPWR VPWR U$$3972/A sky130_fd_sc_hd__buf_4
Xfanout1318 input51/X VGND VGND VPWR VPWR U$$3792/B sky130_fd_sc_hd__buf_6
Xdadda_fa_1_71_0 U$$2144/X U$$2277/X U$$2410/X VGND VGND VPWR VPWR dadda_fa_2_72_0/B
+ dadda_fa_2_71_3/B sky130_fd_sc_hd__fa_1
Xfanout1329 U$$3607/B VGND VGND VPWR VPWR U$$3641/B sky130_fd_sc_hd__buf_6
XFILLER_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout386 U$$1075/A2 VGND VGND VPWR VPWR U$$999/A2 sky130_fd_sc_hd__buf_6
XFILLER_101_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout397 U$$952/A2 VGND VGND VPWR VPWR U$$904/A2 sky130_fd_sc_hd__buf_4
XU$$3109 U$$3109/A U$$3151/A VGND VGND VPWR VPWR U$$3109/X sky130_fd_sc_hd__xor2_1
XFILLER_86_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2408 U$$2408/A U$$2408/B VGND VGND VPWR VPWR U$$2408/X sky130_fd_sc_hd__xor2_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2419 U$$4198/B1 U$$2459/A2 U$$4476/A1 U$$2459/B2 VGND VGND VPWR VPWR U$$2420/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1707 U$$1707/A U$$1721/B VGND VGND VPWR VPWR U$$1707/X sky130_fd_sc_hd__xor2_1
XFILLER_43_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1718 U$$2814/A1 U$$1720/A2 U$$74/B1 U$$1720/B2 VGND VGND VPWR VPWR U$$1719/A sky130_fd_sc_hd__a22o_1
XU$$1729 U$$1729/A U$$1741/B VGND VGND VPWR VPWR U$$1729/X sky130_fd_sc_hd__xor2_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_313_ _321_/CLK _313_/D VGND VGND VPWR VPWR _313_/Q sky130_fd_sc_hd__dfxtp_1
XU$$4461_1878 VGND VGND VPWR VPWR U$$4461_1878/HI U$$4461/B sky130_fd_sc_hd__conb_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_244_ _375_/CLK _244_/D VGND VGND VPWR VPWR _244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput17 a[24] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 a[34] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
Xinput39 a[44] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__dlymetal6s2s_1
X_175_ _319_/CLK _175_/D VGND VGND VPWR VPWR _175_/Q sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_3_93_1 dadda_fa_3_93_1/A dadda_fa_3_93_1/B dadda_fa_3_93_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_0/CIN dadda_fa_4_93_2/A sky130_fd_sc_hd__fa_1
XFILLER_109_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_70_0 dadda_fa_6_70_0/A dadda_fa_6_70_0/B dadda_fa_6_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_71_0/B dadda_fa_7_70_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_86_0 dadda_fa_3_86_0/A dadda_fa_3_86_0/B dadda_fa_3_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_0/B dadda_fa_4_86_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_112_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_2_108_0_1944 VGND VGND VPWR VPWR dadda_ha_2_108_0/A dadda_ha_2_108_0_1944/LO
+ sky130_fd_sc_hd__conb_1
XU$$4300 U$$4300/A U$$4384/A VGND VGND VPWR VPWR U$$4300/X sky130_fd_sc_hd__xor2_1
XFILLER_120_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4311 U$$4446/B1 U$$4373/A2 U$$4450/A1 U$$4373/B2 VGND VGND VPWR VPWR U$$4312/A
+ sky130_fd_sc_hd__a22o_1
XU$$4322 U$$4322/A U$$4322/B VGND VGND VPWR VPWR U$$4322/X sky130_fd_sc_hd__xor2_1
XU$$4333 U$$4470/A1 U$$4349/A2 U$$4472/A1 U$$4349/B2 VGND VGND VPWR VPWR U$$4334/A
+ sky130_fd_sc_hd__a22o_1
XU$$4344 U$$4344/A U$$4350/B VGND VGND VPWR VPWR U$$4344/X sky130_fd_sc_hd__xor2_1
XU$$4355 U$$4492/A1 U$$4359/A2 U$$4492/B1 U$$4359/B2 VGND VGND VPWR VPWR U$$4356/A
+ sky130_fd_sc_hd__a22o_1
XU$$3610 U$$4432/A1 U$$3656/A2 U$$3610/B1 U$$3656/B2 VGND VGND VPWR VPWR U$$3611/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_48_5 dadda_fa_2_48_5/A dadda_fa_2_48_5/B dadda_fa_2_48_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_2/A dadda_fa_4_48_0/A sky130_fd_sc_hd__fa_1
XU$$3621 U$$3621/A U$$3699/A VGND VGND VPWR VPWR U$$3621/X sky130_fd_sc_hd__xor2_1
XFILLER_93_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_115_0 U$$3961/X U$$4094/X U$$4227/X VGND VGND VPWR VPWR dadda_fa_5_116_0/A
+ dadda_fa_5_115_1/A sky130_fd_sc_hd__fa_1
XU$$4366 U$$4366/A U$$4368/B VGND VGND VPWR VPWR U$$4366/X sky130_fd_sc_hd__xor2_1
XU$$3632 U$$4043/A1 U$$3640/A2 U$$4043/B1 U$$3640/B2 VGND VGND VPWR VPWR U$$3633/A
+ sky130_fd_sc_hd__a22o_1
XU$$4377 U$$4512/B1 U$$4381/A2 U$$4377/B1 U$$4381/B2 VGND VGND VPWR VPWR U$$4378/A
+ sky130_fd_sc_hd__a22o_1
XU$$4388 U$$4386/Y U$$4388/A2 U$$4384/A U$$4387/X U$$4384/Y VGND VGND VPWR VPWR U$$4388/X
+ sky130_fd_sc_hd__a32o_1
XU$$3643 U$$3643/A U$$3699/A VGND VGND VPWR VPWR U$$3643/X sky130_fd_sc_hd__xor2_1
XU$$4399 U$$4399/A U$$4399/B VGND VGND VPWR VPWR U$$4399/X sky130_fd_sc_hd__xor2_1
XU$$3654 U$$640/A1 U$$3656/A2 U$$916/A1 U$$3656/B2 VGND VGND VPWR VPWR U$$3655/A sky130_fd_sc_hd__a22o_1
XU$$3665 U$$3665/A U$$3681/B VGND VGND VPWR VPWR U$$3665/X sky130_fd_sc_hd__xor2_1
XU$$2920 U$$2920/A U$$2938/B VGND VGND VPWR VPWR U$$2920/X sky130_fd_sc_hd__xor2_1
XFILLER_34_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2931 U$$4162/B1 U$$2937/A2 U$$4027/B1 U$$2937/B2 VGND VGND VPWR VPWR U$$2932/A
+ sky130_fd_sc_hd__a22o_1
XU$$3676 U$$4359/B1 U$$3692/A2 U$$4226/A1 U$$3692/B2 VGND VGND VPWR VPWR U$$3677/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2942 U$$2942/A U$$2944/B VGND VGND VPWR VPWR U$$2942/X sky130_fd_sc_hd__xor2_1
XU$$3687 U$$3687/A U$$3695/B VGND VGND VPWR VPWR U$$3687/X sky130_fd_sc_hd__xor2_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3698 U$$3698/A VGND VGND VPWR VPWR U$$3698/Y sky130_fd_sc_hd__inv_1
XU$$2953 U$$4049/A1 U$$3005/A2 U$$4460/B1 U$$3005/B2 VGND VGND VPWR VPWR U$$2954/A
+ sky130_fd_sc_hd__a22o_1
XU$$2964 U$$2964/A U$$2974/B VGND VGND VPWR VPWR U$$2964/X sky130_fd_sc_hd__xor2_1
XFILLER_61_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2975 U$$3112/A1 U$$2977/A2 U$$922/A1 U$$2977/B2 VGND VGND VPWR VPWR U$$2976/A
+ sky130_fd_sc_hd__a22o_1
XU$$2986 U$$2986/A U$$2986/B VGND VGND VPWR VPWR U$$2986/X sky130_fd_sc_hd__xor2_1
XFILLER_60_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2997 U$$3817/B1 U$$3005/A2 U$$3684/A1 U$$3005/B2 VGND VGND VPWR VPWR U$$2998/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$915 final_adder.U$$144/A final_adder.U$$853/X final_adder.U$$915/B1
+ VGND VGND VPWR VPWR final_adder.U$$915/X sky130_fd_sc_hd__a21o_1
XFILLER_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$937 final_adder.U$$166/A final_adder.U$$875/X final_adder.U$$937/B1
+ VGND VGND VPWR VPWR final_adder.U$$937/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_5 U$$2102/X U$$2235/X U$$2368/X VGND VGND VPWR VPWR dadda_fa_2_51_2/A
+ dadda_fa_2_50_5/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$959 final_adder.U$$188/A final_adder.U$$897/X final_adder.U$$959/B1
+ VGND VGND VPWR VPWR final_adder.U$$959/X sky130_fd_sc_hd__a21o_1
XU$$809 U$$944/B1 U$$809/A2 U$$811/A1 U$$809/B2 VGND VGND VPWR VPWR U$$810/A sky130_fd_sc_hd__a22o_1
XFILLER_56_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1104 input80/X VGND VGND VPWR VPWR U$$602/A1 sky130_fd_sc_hd__buf_4
Xfanout1115 U$$3751/A1 VGND VGND VPWR VPWR U$$4162/A1 sky130_fd_sc_hd__buf_6
XFILLER_154_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1126 U$$2925/A1 VGND VGND VPWR VPWR U$$596/A1 sky130_fd_sc_hd__buf_4
XFILLER_121_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1137 U$$3846/A1 VGND VGND VPWR VPWR U$$969/A1 sky130_fd_sc_hd__buf_4
Xfanout1148 U$$4017/B1 VGND VGND VPWR VPWR U$$183/A1 sky130_fd_sc_hd__buf_4
Xfanout1159 U$$3056/A1 VGND VGND VPWR VPWR U$$864/A1 sky130_fd_sc_hd__buf_4
XFILLER_59_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2205 U$$2205/A U$$2253/B VGND VGND VPWR VPWR U$$2205/X sky130_fd_sc_hd__xor2_1
XFILLER_90_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2216 U$$983/A1 U$$2254/A2 U$$983/B1 U$$2254/B2 VGND VGND VPWR VPWR U$$2217/A sky130_fd_sc_hd__a22o_1
XU$$2227 U$$2227/A U$$2231/B VGND VGND VPWR VPWR U$$2227/X sky130_fd_sc_hd__xor2_1
XFILLER_28_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2238 U$$183/A1 U$$2248/A2 U$$870/A1 U$$2248/B2 VGND VGND VPWR VPWR U$$2239/A sky130_fd_sc_hd__a22o_1
XU$$1504 U$$4244/A1 U$$1504/A2 U$$1504/B1 U$$1504/B2 VGND VGND VPWR VPWR U$$1505/A
+ sky130_fd_sc_hd__a22o_1
XU$$2249 U$$2249/A U$$2249/B VGND VGND VPWR VPWR U$$2249/X sky130_fd_sc_hd__xor2_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1515 U$$2748/A1 U$$1575/A2 U$$3296/B1 U$$1575/B2 VGND VGND VPWR VPWR U$$1516/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1526 U$$1526/A U$$1564/B VGND VGND VPWR VPWR U$$1526/X sky130_fd_sc_hd__xor2_1
XFILLER_15_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1537 U$$30/A1 U$$1575/A2 U$$32/A1 U$$1575/B2 VGND VGND VPWR VPWR U$$1538/A sky130_fd_sc_hd__a22o_1
XU$$1548 U$$1548/A U$$1570/B VGND VGND VPWR VPWR U$$1548/X sky130_fd_sc_hd__xor2_1
XU$$1559 U$$598/B1 U$$1563/A2 U$$465/A1 U$$1563/B2 VGND VGND VPWR VPWR U$$1560/A sky130_fd_sc_hd__a22o_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_227_ _356_/CLK _227_/D VGND VGND VPWR VPWR _227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_60_4 dadda_fa_2_60_4/A dadda_fa_2_60_4/B dadda_fa_2_60_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_1/CIN dadda_fa_3_60_3/CIN sky130_fd_sc_hd__fa_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1660 U$$4496/A1 VGND VGND VPWR VPWR U$$3948/A1 sky130_fd_sc_hd__buf_4
XFILLER_38_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_53_3 dadda_fa_2_53_3/A dadda_fa_2_53_3/B dadda_fa_2_53_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_1/B dadda_fa_3_53_3/B sky130_fd_sc_hd__fa_1
Xfanout1671 U$$2711/B1 VGND VGND VPWR VPWR U$$4494/A1 sky130_fd_sc_hd__buf_4
Xfanout1682 U$$1328/B VGND VGND VPWR VPWR U$$1294/B sky130_fd_sc_hd__clkbuf_8
XU$$4130 U$$4265/B1 U$$4158/A2 U$$4132/A1 U$$4158/B2 VGND VGND VPWR VPWR U$$4131/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1693 U$$3850/B1 VGND VGND VPWR VPWR U$$3030/A1 sky130_fd_sc_hd__buf_4
XU$$4141 U$$4141/A U$$4191/B VGND VGND VPWR VPWR U$$4141/X sky130_fd_sc_hd__xor2_1
XU$$4152 U$$4152/A1 U$$4244/A2 U$$4152/B1 U$$4244/B2 VGND VGND VPWR VPWR U$$4153/A
+ sky130_fd_sc_hd__a22o_1
XU$$4163 U$$4163/A U$$4175/B VGND VGND VPWR VPWR U$$4163/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_46_2 dadda_fa_2_46_2/A dadda_fa_2_46_2/B dadda_fa_2_46_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_1/A dadda_fa_3_46_3/A sky130_fd_sc_hd__fa_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4174 U$$4174/A1 U$$4174/A2 U$$4176/A1 U$$4174/B2 VGND VGND VPWR VPWR U$$4175/A
+ sky130_fd_sc_hd__a22o_1
XU$$3440 U$$3440/A U$$3482/B VGND VGND VPWR VPWR U$$3440/X sky130_fd_sc_hd__xor2_1
XFILLER_168_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_23_1 dadda_fa_5_23_1/A dadda_fa_5_23_1/B dadda_fa_5_23_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_24_0/B dadda_fa_7_23_0/A sky130_fd_sc_hd__fa_2
XU$$4185 U$$4185/A U$$4215/B VGND VGND VPWR VPWR U$$4185/X sky130_fd_sc_hd__xor2_1
XU$$3451 U$$3999/A1 U$$3473/A2 U$$3999/B1 U$$3473/B2 VGND VGND VPWR VPWR U$$3452/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_39_1 U$$1548/X U$$1681/X U$$1814/X VGND VGND VPWR VPWR dadda_fa_3_40_0/CIN
+ dadda_fa_3_39_2/CIN sky130_fd_sc_hd__fa_1
XU$$4196 U$$4196/A1 U$$4224/A2 U$$4196/B1 U$$4224/B2 VGND VGND VPWR VPWR U$$4197/A
+ sky130_fd_sc_hd__a22o_1
XU$$3462 U$$3462/A U$$3468/B VGND VGND VPWR VPWR U$$3462/X sky130_fd_sc_hd__xor2_1
XU$$3473 U$$4432/A1 U$$3473/A2 U$$872/A1 U$$3473/B2 VGND VGND VPWR VPWR U$$3474/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3484 U$$3484/A U$$3558/B VGND VGND VPWR VPWR U$$3484/X sky130_fd_sc_hd__xor2_1
XU$$2750 U$$3022/B1 U$$2798/A2 U$$2887/B1 U$$2798/B2 VGND VGND VPWR VPWR U$$2751/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_16_0 dadda_fa_5_16_0/A dadda_fa_5_16_0/B dadda_fa_5_16_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_17_0/A dadda_fa_6_16_0/CIN sky130_fd_sc_hd__fa_1
XU$$3495 U$$3630/B1 U$$3505/A2 U$$3495/B1 U$$3505/B2 VGND VGND VPWR VPWR U$$3496/A
+ sky130_fd_sc_hd__a22o_1
XU$$2761 U$$2761/A U$$2799/B VGND VGND VPWR VPWR U$$2761/X sky130_fd_sc_hd__xor2_1
XU$$2772 U$$32/A1 U$$2812/A2 U$$32/B1 U$$2812/B2 VGND VGND VPWR VPWR U$$2773/A sky130_fd_sc_hd__a22o_1
XU$$2783 U$$2783/A U$$2811/B VGND VGND VPWR VPWR U$$2783/X sky130_fd_sc_hd__xor2_1
XU$$2794 U$$602/A1 U$$2798/A2 U$$3205/B1 U$$2798/B2 VGND VGND VPWR VPWR U$$2795/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput207 c[55] VGND VGND VPWR VPWR input207/X sky130_fd_sc_hd__clkbuf_4
Xinput218 c[65] VGND VGND VPWR VPWR input218/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput229 c[75] VGND VGND VPWR VPWR input229/X sky130_fd_sc_hd__buf_2
Xfinal_adder.U$$701 final_adder.U$$700/B final_adder.U$$597/X final_adder.U$$581/X
+ VGND VGND VPWR VPWR final_adder.U$$701/X sky130_fd_sc_hd__a21o_1
XFILLER_124_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$712 final_adder.U$$712/A final_adder.U$$712/B VGND VGND VPWR VPWR
+ final_adder.U$$792/A sky130_fd_sc_hd__and2_1
XFILLER_97_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$723 final_adder.U$$706/A final_adder.U$$619/X final_adder.U$$603/X
+ VGND VGND VPWR VPWR final_adder.U$$723/X sky130_fd_sc_hd__a21o_2
XFILLER_112_1012 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$745 final_adder.U$$744/B final_adder.U$$665/X final_adder.U$$633/X
+ VGND VGND VPWR VPWR final_adder.U$$745/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$756 final_adder.U$$788/B final_adder.U$$756/B VGND VGND VPWR VPWR
+ final_adder.U$$756/X sky130_fd_sc_hd__and2_1
XFILLER_57_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$767 final_adder.U$$766/B final_adder.U$$687/X final_adder.U$$655/X
+ VGND VGND VPWR VPWR final_adder.U$$767/X sky130_fd_sc_hd__a21o_1
XU$$606 U$$880/A1 U$$638/A2 U$$882/A1 U$$638/B2 VGND VGND VPWR VPWR U$$607/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$778 final_adder.U$$778/A final_adder.U$$778/B VGND VGND VPWR VPWR
+ final_adder.U$$778/X sky130_fd_sc_hd__and2_1
XFILLER_44_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$617 U$$617/A U$$637/B VGND VGND VPWR VPWR U$$617/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$789 final_adder.U$$788/B final_adder.U$$709/X final_adder.U$$677/X
+ VGND VGND VPWR VPWR final_adder.U$$789/X sky130_fd_sc_hd__a21o_1
XU$$628 U$$900/B1 U$$630/A2 U$$765/B1 U$$630/B2 VGND VGND VPWR VPWR U$$629/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_41_1 U$$488/X U$$621/X U$$754/X VGND VGND VPWR VPWR dadda_fa_2_42_3/CIN
+ dadda_fa_2_41_5/B sky130_fd_sc_hd__fa_1
XFILLER_72_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$639 U$$639/A U$$639/B VGND VGND VPWR VPWR U$$639/X sky130_fd_sc_hd__xor2_1
XFILLER_83_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1915_1795 VGND VGND VPWR VPWR U$$1915_1795/HI U$$1915/B1 sky130_fd_sc_hd__conb_1
XFILLER_138_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_70_3 dadda_fa_3_70_3/A dadda_fa_3_70_3/B dadda_fa_3_70_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_1/B dadda_fa_4_70_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_63_2 dadda_fa_3_63_2/A dadda_fa_3_63_2/B dadda_fa_3_63_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_1/A dadda_fa_4_63_2/B sky130_fd_sc_hd__fa_1
XFILLER_0_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_56_1 dadda_fa_3_56_1/A dadda_fa_3_56_1/B dadda_fa_3_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_0/CIN dadda_fa_4_56_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_33_0 dadda_fa_6_33_0/A dadda_fa_6_33_0/B dadda_fa_6_33_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_34_0/B dadda_fa_7_33_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_49_0 dadda_fa_3_49_0/A dadda_fa_3_49_0/B dadda_fa_3_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_0/B dadda_fa_4_49_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2002 U$$3509/A1 U$$2046/A2 U$$86/A1 U$$2046/B2 VGND VGND VPWR VPWR U$$2003/A sky130_fd_sc_hd__a22o_1
XU$$2013 U$$2013/A U$$2015/B VGND VGND VPWR VPWR U$$2013/X sky130_fd_sc_hd__xor2_1
XU$$2024 U$$4353/A1 U$$2052/A2 U$$4353/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2025/A
+ sky130_fd_sc_hd__a22o_1
XU$$2035 U$$2035/A U$$2043/B VGND VGND VPWR VPWR U$$2035/X sky130_fd_sc_hd__xor2_1
XFILLER_63_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1301 U$$66/B1 U$$1327/A2 U$$892/A1 U$$1327/B2 VGND VGND VPWR VPWR U$$1302/A sky130_fd_sc_hd__a22o_1
XU$$2046 U$$2183/A1 U$$2046/A2 U$$4512/B1 U$$2046/B2 VGND VGND VPWR VPWR U$$2047/A
+ sky130_fd_sc_hd__a22o_1
XU$$2057 U$$2192/A VGND VGND VPWR VPWR U$$2057/Y sky130_fd_sc_hd__inv_1
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1312 U$$1312/A U$$1320/B VGND VGND VPWR VPWR U$$1312/X sky130_fd_sc_hd__xor2_1
XU$$1323 U$$90/A1 U$$1367/A2 U$$92/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1324/A sky130_fd_sc_hd__a22o_1
XU$$2068 U$$2068/A U$$2106/B VGND VGND VPWR VPWR U$$2068/X sky130_fd_sc_hd__xor2_1
XU$$1334 U$$1334/A U$$1370/A VGND VGND VPWR VPWR U$$1334/X sky130_fd_sc_hd__xor2_1
XU$$2079 U$$981/B1 U$$2107/A2 U$$2629/A1 U$$2107/B2 VGND VGND VPWR VPWR U$$2080/A
+ sky130_fd_sc_hd__a22o_1
XU$$1345 U$$521/B1 U$$1359/A2 U$$386/B1 U$$1359/B2 VGND VGND VPWR VPWR U$$1346/A sky130_fd_sc_hd__a22o_1
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1356 U$$1356/A U$$1358/B VGND VGND VPWR VPWR U$$1356/X sky130_fd_sc_hd__xor2_1
XU$$1367 U$$406/B1 U$$1367/A2 U$$1367/B1 U$$1367/B2 VGND VGND VPWR VPWR U$$1368/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_114_1 U$$3826/X U$$3959/X VGND VGND VPWR VPWR dadda_fa_4_115_2/B dadda_ha_3_114_1/SUM
+ sky130_fd_sc_hd__ha_1
XU$$1378 U$$828/B1 U$$1414/A2 U$$3435/A1 U$$1414/B2 VGND VGND VPWR VPWR U$$1379/A
+ sky130_fd_sc_hd__a22o_1
XU$$1389 U$$1389/A U$$1427/B VGND VGND VPWR VPWR U$$1389/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_106_0 dadda_fa_7_106_0/A dadda_fa_7_106_0/B dadda_fa_7_106_0/CIN VGND
+ VGND VPWR VPWR _403_/D _274_/D sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_10_clk _201_/CLK VGND VGND VPWR VPWR _359_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1150 final_adder.U$$899/A1 final_adder.U$$837/X VGND VGND VPWR VPWR
+ output286/A sky130_fd_sc_hd__xor2_4
XFILLER_116_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout908 U$$1218/B2 VGND VGND VPWR VPWR U$$1170/B2 sky130_fd_sc_hd__buf_4
XFILLER_124_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout919 U$$102/B2 VGND VGND VPWR VPWR U$$120/B2 sky130_fd_sc_hd__buf_6
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_51_0 input203/X dadda_fa_2_51_0/B dadda_fa_2_51_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_52_0/B dadda_fa_3_51_2/B sky130_fd_sc_hd__fa_1
Xfanout1490 U$$1618/B VGND VGND VPWR VPWR U$$1584/B sky130_fd_sc_hd__buf_6
XFILLER_54_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$30 _326_/Q _198_/Q VGND VGND VPWR VPWR final_adder.U$$995/B1 final_adder.U$$224/A
+ sky130_fd_sc_hd__ha_1
XFILLER_80_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$41 _337_/Q _209_/Q VGND VGND VPWR VPWR final_adder.U$$215/B1 final_adder.U$$214/B
+ sky130_fd_sc_hd__ha_1
XFILLER_54_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3270 U$$3270/A U$$3286/B VGND VGND VPWR VPWR U$$3270/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$52 _348_/Q _220_/Q VGND VGND VPWR VPWR final_adder.U$$973/B1 final_adder.U$$202/A
+ sky130_fd_sc_hd__ha_2
XFILLER_0_1044 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3281 U$$3418/A1 U$$3283/A2 U$$3418/B1 U$$3283/B2 VGND VGND VPWR VPWR U$$3282/A
+ sky130_fd_sc_hd__a22o_1
XU$$3292 U$$3290/Y input43/X U$$3288/A U$$3291/X U$$3288/Y VGND VGND VPWR VPWR U$$3292/X
+ sky130_fd_sc_hd__a32o_4
Xfinal_adder.U$$63 _359_/Q _231_/Q VGND VGND VPWR VPWR final_adder.U$$193/B1 final_adder.U$$192/B
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$74 _370_/Q _242_/Q VGND VGND VPWR VPWR final_adder.U$$951/B1 final_adder.U$$180/A
+ sky130_fd_sc_hd__ha_1
XFILLER_94_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$85 _381_/Q _253_/Q VGND VGND VPWR VPWR final_adder.U$$171/B1 final_adder.U$$170/B
+ sky130_fd_sc_hd__ha_2
XFILLER_81_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$96 _392_/Q _264_/Q VGND VGND VPWR VPWR final_adder.U$$929/B1 final_adder.U$$158/A
+ sky130_fd_sc_hd__ha_1
XU$$2580 U$$4361/A1 U$$2598/A2 U$$4363/A1 U$$2598/B2 VGND VGND VPWR VPWR U$$2581/A
+ sky130_fd_sc_hd__a22o_1
XU$$2591 U$$2591/A U$$2591/B VGND VGND VPWR VPWR U$$2591/X sky130_fd_sc_hd__xor2_1
XFILLER_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1890 U$$1890/A U$$1916/B VGND VGND VPWR VPWR U$$1890/X sky130_fd_sc_hd__xor2_1
XFILLER_119_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_80_2 dadda_fa_4_80_2/A dadda_fa_4_80_2/B dadda_fa_4_80_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_81_0/CIN dadda_fa_5_80_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_73_1 dadda_fa_4_73_1/A dadda_fa_4_73_1/B dadda_fa_4_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_74_0/B dadda_fa_5_73_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_89_1 U$$2180/X U$$2313/X U$$2446/X VGND VGND VPWR VPWR dadda_fa_2_90_4/A
+ dadda_fa_2_89_5/B sky130_fd_sc_hd__fa_1
XFILLER_116_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_50_0 dadda_fa_7_50_0/A dadda_fa_7_50_0/B dadda_fa_7_50_0/CIN VGND VGND
+ VPWR VPWR _347_/D _218_/D sky130_fd_sc_hd__fa_2
XFILLER_135_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_66_0 dadda_fa_4_66_0/A dadda_fa_4_66_0/B dadda_fa_4_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_67_0/A dadda_fa_5_66_1/A sky130_fd_sc_hd__fa_1
XFILLER_131_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$520 final_adder.U$$528/B final_adder.U$$520/B VGND VGND VPWR VPWR
+ final_adder.U$$640/B sky130_fd_sc_hd__and2_1
XFILLER_85_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$531 final_adder.U$$530/B final_adder.U$$415/X final_adder.U$$407/X
+ VGND VGND VPWR VPWR final_adder.U$$531/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$542 final_adder.U$$550/B final_adder.U$$542/B VGND VGND VPWR VPWR
+ final_adder.U$$662/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$553 final_adder.U$$552/B final_adder.U$$437/X final_adder.U$$429/X
+ VGND VGND VPWR VPWR final_adder.U$$553/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$564 final_adder.U$$572/B final_adder.U$$564/B VGND VGND VPWR VPWR
+ final_adder.U$$684/B sky130_fd_sc_hd__and2_1
XU$$403 U$$403/A U$$411/A VGND VGND VPWR VPWR U$$403/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$575 final_adder.U$$574/B final_adder.U$$459/X final_adder.U$$451/X
+ VGND VGND VPWR VPWR final_adder.U$$575/X sky130_fd_sc_hd__a21o_1
XU$$414 U$$536/B U$$414/B VGND VGND VPWR VPWR U$$414/X sky130_fd_sc_hd__and2_1
XFILLER_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$586 final_adder.U$$594/B final_adder.U$$586/B VGND VGND VPWR VPWR
+ final_adder.U$$706/B sky130_fd_sc_hd__and2_1
XU$$425 U$$14/A1 U$$479/A2 U$$16/A1 U$$479/B2 VGND VGND VPWR VPWR U$$426/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$597 final_adder.U$$596/B final_adder.U$$481/X final_adder.U$$473/X
+ VGND VGND VPWR VPWR final_adder.U$$597/X sky130_fd_sc_hd__a21o_1
XU$$436 U$$436/A U$$506/B VGND VGND VPWR VPWR U$$436/X sky130_fd_sc_hd__xor2_1
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$447 U$$447/A1 U$$447/A2 U$$447/B1 U$$447/B2 VGND VGND VPWR VPWR U$$448/A sky130_fd_sc_hd__a22o_1
XU$$458 U$$458/A U$$498/B VGND VGND VPWR VPWR U$$458/X sky130_fd_sc_hd__xor2_1
XFILLER_60_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$469 U$$56/B1 U$$501/A2 U$$469/B1 U$$501/B2 VGND VGND VPWR VPWR U$$470/A sky130_fd_sc_hd__a22o_1
XFILLER_71_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$970 U$$970/A U$$982/B VGND VGND VPWR VPWR U$$970/X sky130_fd_sc_hd__xor2_1
XU$$1120 U$$981/B1 U$$1194/A2 U$$2629/A1 U$$1194/B2 VGND VGND VPWR VPWR U$$1121/A
+ sky130_fd_sc_hd__a22o_1
XU$$981 U$$981/A1 U$$981/A2 U$$981/B1 U$$981/B2 VGND VGND VPWR VPWR U$$982/A sky130_fd_sc_hd__a22o_1
XU$$992 U$$992/A U$$998/B VGND VGND VPWR VPWR U$$992/X sky130_fd_sc_hd__xor2_1
XU$$1131 U$$1131/A U$$1163/B VGND VGND VPWR VPWR U$$1131/X sky130_fd_sc_hd__xor2_1
XFILLER_90_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1142 U$$46/A1 U$$1174/A2 U$$48/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1143/A sky130_fd_sc_hd__a22o_1
XU$$1153 U$$1153/A U$$1195/B VGND VGND VPWR VPWR U$$1153/X sky130_fd_sc_hd__xor2_1
XU$$1164 U$$66/B1 U$$1164/A2 U$$892/A1 U$$1164/B2 VGND VGND VPWR VPWR U$$1165/A sky130_fd_sc_hd__a22o_1
XU$$3157_1816 VGND VGND VPWR VPWR U$$3157_1816/HI U$$3157/A1 sky130_fd_sc_hd__conb_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1175 U$$1175/A U$$1175/B VGND VGND VPWR VPWR U$$1175/X sky130_fd_sc_hd__xor2_1
XU$$1186 U$$773/B1 U$$1226/A2 U$$640/A1 U$$1226/B2 VGND VGND VPWR VPWR U$$1187/A sky130_fd_sc_hd__a22o_1
XFILLER_148_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1197 U$$1197/A U$$1233/A VGND VGND VPWR VPWR U$$1197/X sky130_fd_sc_hd__xor2_1
XFILLER_129_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_90_1 dadda_fa_5_90_1/A dadda_fa_5_90_1/B dadda_fa_5_90_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_91_0/B dadda_fa_7_90_0/A sky130_fd_sc_hd__fa_1
XFILLER_117_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_83_0 dadda_fa_5_83_0/A dadda_fa_5_83_0/B dadda_fa_5_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_84_0/A dadda_fa_6_83_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_99_0 U$$2465/Y U$$2599/X U$$2732/X VGND VGND VPWR VPWR dadda_fa_3_100_1/A
+ dadda_fa_3_99_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout705 U$$4115/X VGND VGND VPWR VPWR U$$4236/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout716 U$$4057/B2 VGND VGND VPWR VPWR U$$4093/B2 sky130_fd_sc_hd__buf_2
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout727 U$$3777/B2 VGND VGND VPWR VPWR U$$3757/B2 sky130_fd_sc_hd__buf_4
XFILLER_59_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_75_7 U$$4413/X input229/X dadda_fa_1_75_7/CIN VGND VGND VPWR VPWR dadda_fa_2_76_2/CIN
+ dadda_fa_2_75_5/CIN sky130_fd_sc_hd__fa_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout738 U$$3658/B2 VGND VGND VPWR VPWR U$$3656/B2 sky130_fd_sc_hd__buf_4
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 U$$3557/B2 VGND VGND VPWR VPWR U$$3559/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_6 dadda_fa_1_68_6/A dadda_fa_1_68_6/B dadda_fa_1_68_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_69_2/B dadda_fa_2_68_5/B sky130_fd_sc_hd__fa_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_942 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_98_0 dadda_fa_7_98_0/A dadda_fa_7_98_0/B dadda_fa_7_98_0/CIN VGND VGND
+ VPWR VPWR _395_/D _266_/D sky130_fd_sc_hd__fa_1
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_113_0 dadda_fa_6_113_0/A dadda_fa_6_113_0/B dadda_fa_6_113_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_114_0/B dadda_fa_7_113_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$350 final_adder.U$$352/B final_adder.U$$350/B VGND VGND VPWR VPWR
+ final_adder.U$$476/B sky130_fd_sc_hd__and2_1
XFILLER_92_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$361 final_adder.U$$360/B final_adder.U$$235/X final_adder.U$$233/X
+ VGND VGND VPWR VPWR final_adder.U$$361/X sky130_fd_sc_hd__a21o_1
XU$$200 U$$200/A U$$230/B VGND VGND VPWR VPWR U$$200/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$372 final_adder.U$$374/B final_adder.U$$372/B VGND VGND VPWR VPWR
+ final_adder.U$$498/B sky130_fd_sc_hd__and2_1
XU$$211 U$$74/A1 U$$213/A2 U$$76/A1 U$$213/B2 VGND VGND VPWR VPWR U$$212/A sky130_fd_sc_hd__a22o_1
XU$$222 U$$222/A U$$230/B VGND VGND VPWR VPWR U$$222/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_33_3 dadda_fa_3_33_3/A dadda_fa_3_33_3/B dadda_fa_3_33_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_34_1/B dadda_fa_4_33_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$394 final_adder.U$$398/B final_adder.U$$394/B VGND VGND VPWR VPWR
+ final_adder.U$$518/B sky130_fd_sc_hd__and2_1
XU$$233 U$$96/A1 U$$271/A2 U$$98/A1 U$$271/B2 VGND VGND VPWR VPWR U$$234/A sky130_fd_sc_hd__a22o_1
XFILLER_73_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$244 U$$244/A U$$254/B VGND VGND VPWR VPWR U$$244/X sky130_fd_sc_hd__xor2_1
XU$$255 U$$803/A1 U$$259/A2 U$$942/A1 U$$259/B2 VGND VGND VPWR VPWR U$$256/A sky130_fd_sc_hd__a22o_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_26_2 U$$1828/B input175/X dadda_fa_3_26_2/CIN VGND VGND VPWR VPWR dadda_fa_4_27_1/A
+ dadda_fa_4_26_2/B sky130_fd_sc_hd__fa_1
XU$$266 U$$266/A U$$274/A VGND VGND VPWR VPWR U$$266/X sky130_fd_sc_hd__xor2_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$277 U$$411/A U$$277/B VGND VGND VPWR VPWR U$$277/X sky130_fd_sc_hd__and2_1
XFILLER_72_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$288 U$$14/A1 U$$312/A2 U$$16/A1 U$$312/B2 VGND VGND VPWR VPWR U$$289/A sky130_fd_sc_hd__a22o_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_19_1 U$$444/X U$$577/X U$$710/X VGND VGND VPWR VPWR dadda_fa_4_20_1/A
+ dadda_fa_4_19_2/B sky130_fd_sc_hd__fa_1
XU$$299 U$$299/A U$$341/B VGND VGND VPWR VPWR U$$299/X sky130_fd_sc_hd__xor2_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$5 U$$3/B U$$5/A2 U$$1/A U$$0/Y VGND VGND VPWR VPWR U$$5/X sky130_fd_sc_hd__a22o_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput308 output308/A VGND VGND VPWR VPWR o[30] sky130_fd_sc_hd__buf_2
Xoutput319 output319/A VGND VGND VPWR VPWR o[40] sky130_fd_sc_hd__buf_2
XFILLER_114_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_78_5 dadda_fa_2_78_5/A dadda_fa_2_78_5/B dadda_fa_2_78_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_2/A dadda_fa_4_78_0/A sky130_fd_sc_hd__fa_2
XFILLER_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_839 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_108_1 dadda_fa_5_108_1/A dadda_fa_5_108_1/B dadda_fa_5_108_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_109_0/B dadda_fa_7_108_0/A sky130_fd_sc_hd__fa_1
XFILLER_117_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_80_5 U$$3093/X U$$3226/X U$$3359/X VGND VGND VPWR VPWR dadda_fa_2_81_2/B
+ dadda_fa_2_80_5/A sky130_fd_sc_hd__fa_1
XFILLER_104_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout502 U$$3207/A2 VGND VGND VPWR VPWR U$$3199/A2 sky130_fd_sc_hd__buf_6
Xfanout513 U$$3112/A2 VGND VGND VPWR VPWR U$$3108/A2 sky130_fd_sc_hd__buf_4
Xfanout524 U$$2881/X VGND VGND VPWR VPWR U$$2991/A2 sky130_fd_sc_hd__buf_6
XFILLER_116_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_73_4 U$$3478/X U$$3611/X U$$3744/X VGND VGND VPWR VPWR dadda_fa_2_74_1/CIN
+ dadda_fa_2_73_4/CIN sky130_fd_sc_hd__fa_1
Xfanout535 U$$386/A2 VGND VGND VPWR VPWR U$$338/A2 sky130_fd_sc_hd__buf_2
Xfanout546 U$$2607/X VGND VGND VPWR VPWR U$$2667/A2 sky130_fd_sc_hd__buf_4
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout557 fanout561/X VGND VGND VPWR VPWR U$$2546/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_66_3 U$$3730/X U$$3863/X U$$3996/X VGND VGND VPWR VPWR dadda_fa_2_67_1/B
+ dadda_fa_2_66_4/B sky130_fd_sc_hd__fa_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout568 U$$2463/A2 VGND VGND VPWR VPWR U$$2459/A2 sky130_fd_sc_hd__buf_6
Xfanout579 U$$2059/X VGND VGND VPWR VPWR U$$2139/A2 sky130_fd_sc_hd__clkbuf_8
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_43_2 dadda_fa_4_43_2/A dadda_fa_4_43_2/B dadda_fa_4_43_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_44_0/CIN dadda_fa_5_43_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_59_2 U$$2386/X U$$2519/X U$$2652/X VGND VGND VPWR VPWR dadda_fa_2_60_1/A
+ dadda_fa_2_59_4/A sky130_fd_sc_hd__fa_1
XFILLER_27_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_36_1 dadda_fa_4_36_1/A dadda_fa_4_36_1/B dadda_fa_4_36_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_37_0/B dadda_fa_5_36_1/B sky130_fd_sc_hd__fa_1
XFILLER_27_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_13_0 dadda_fa_7_13_0/A dadda_fa_7_13_0/B dadda_fa_7_13_0/CIN VGND VGND
+ VPWR VPWR _310_/D _181_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_29_0 dadda_fa_4_29_0/A dadda_fa_4_29_0/B dadda_fa_4_29_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_30_0/A dadda_fa_5_29_1/A sky130_fd_sc_hd__fa_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ _391_/CLK _260_/D VGND VGND VPWR VPWR _260_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_191_ _321_/CLK _191_/D VGND VGND VPWR VPWR _191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4504 U$$4504/A1 U$$4388/X U$$4506/A1 U$$4506/B2 VGND VGND VPWR VPWR U$$4505/A
+ sky130_fd_sc_hd__a22o_1
XU$$4515 U$$4515/A U$$4515/B VGND VGND VPWR VPWR U$$4515/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_61_2 U$$927/X U$$1060/X U$$1193/X VGND VGND VPWR VPWR dadda_fa_1_62_6/B
+ dadda_fa_1_61_8/B sky130_fd_sc_hd__fa_1
XU$$3803 U$$4488/A1 U$$3833/A2 U$$4490/A1 U$$3833/B2 VGND VGND VPWR VPWR U$$3804/A
+ sky130_fd_sc_hd__a22o_1
XU$$3814 U$$3814/A U$$3816/B VGND VGND VPWR VPWR U$$3814/X sky130_fd_sc_hd__xor2_1
XU$$18 U$$18/A1 U$$8/A2 U$$20/A1 U$$8/B2 VGND VGND VPWR VPWR U$$19/A sky130_fd_sc_hd__a22o_1
XU$$29 U$$29/A U$$81/B VGND VGND VPWR VPWR U$$29/X sky130_fd_sc_hd__xor2_1
XU$$3825 U$$3960/B1 U$$3825/A2 U$$3825/B1 U$$3825/B2 VGND VGND VPWR VPWR U$$3826/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3836 U$$3836/A VGND VGND VPWR VPWR U$$3836/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_3_31_0 U$$1931/X U$$2064/X input181/X VGND VGND VPWR VPWR dadda_fa_4_32_0/B
+ dadda_fa_4_31_1/CIN sky130_fd_sc_hd__fa_1
XU$$3847 U$$3847/A U$$3893/B VGND VGND VPWR VPWR U$$3847/X sky130_fd_sc_hd__xor2_1
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$180 final_adder.U$$180/A final_adder.U$$180/B VGND VGND VPWR VPWR
+ final_adder.U$$308/B sky130_fd_sc_hd__and2_1
XU$$3858 U$$4132/A1 U$$3892/A2 U$$4132/B1 U$$3892/B2 VGND VGND VPWR VPWR U$$3859/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$191 final_adder.U$$190/B final_adder.U$$961/B1 final_adder.U$$191/B1
+ VGND VGND VPWR VPWR final_adder.U$$191/X sky130_fd_sc_hd__a21o_1
XU$$3869 U$$3869/A U$$3893/B VGND VGND VPWR VPWR U$$3869/X sky130_fd_sc_hd__xor2_1
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_389_ _391_/CLK _389_/D VGND VGND VPWR VPWR _389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_90_4 dadda_fa_2_90_4/A dadda_fa_2_90_4/B dadda_fa_2_90_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_91_1/CIN dadda_fa_3_90_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_127_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_83_3 dadda_fa_2_83_3/A dadda_fa_2_83_3/B dadda_fa_2_83_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_1/B dadda_fa_3_83_3/B sky130_fd_sc_hd__fa_1
XFILLER_88_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_76_2 dadda_fa_2_76_2/A dadda_fa_2_76_2/B dadda_fa_2_76_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_1/A dadda_fa_3_76_3/A sky130_fd_sc_hd__fa_1
XFILLER_87_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_53_1 dadda_fa_5_53_1/A dadda_fa_5_53_1/B dadda_fa_5_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_54_0/B dadda_fa_7_53_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_69_1 dadda_fa_2_69_1/A dadda_fa_2_69_1/B dadda_fa_2_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_0/CIN dadda_fa_3_69_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_46_0 dadda_fa_5_46_0/A dadda_fa_5_46_0/B dadda_fa_5_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_47_0/A dadda_fa_6_46_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4447_1871 VGND VGND VPWR VPWR U$$4447_1871/HI U$$4447/B sky130_fd_sc_hd__conb_1
XFILLER_102_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_120_0 U$$4503/X input152/X dadda_fa_5_120_0/CIN VGND VGND VPWR VPWR dadda_fa_6_121_0/A
+ dadda_fa_6_120_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_104_0_1933 VGND VGND VPWR VPWR dadda_fa_2_104_0/A dadda_fa_2_104_0_1933/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_774 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1308 fanout1309/X VGND VGND VPWR VPWR U$$3925/B sky130_fd_sc_hd__buf_6
Xfanout1319 U$$925/B VGND VGND VPWR VPWR U$$895/B sky130_fd_sc_hd__buf_6
Xdadda_fa_1_71_1 U$$2543/X U$$2676/X U$$2809/X VGND VGND VPWR VPWR dadda_fa_2_72_0/CIN
+ dadda_fa_2_71_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_64_0 U$$2529/X U$$2662/X U$$2795/X VGND VGND VPWR VPWR dadda_fa_2_65_0/B
+ dadda_fa_2_64_3/B sky130_fd_sc_hd__fa_1
Xfanout387 U$$963/X VGND VGND VPWR VPWR U$$1075/A2 sky130_fd_sc_hd__buf_6
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout398 U$$952/A2 VGND VGND VPWR VPWR U$$956/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2409 U$$3916/A1 U$$2459/A2 U$$4466/A1 U$$2459/B2 VGND VGND VPWR VPWR U$$2410/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1708 U$$747/B1 U$$1720/A2 U$$749/B1 U$$1720/B2 VGND VGND VPWR VPWR U$$1709/A sky130_fd_sc_hd__a22o_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1719 U$$1719/A U$$1721/B VGND VGND VPWR VPWR U$$1719/X sky130_fd_sc_hd__xor2_1
XFILLER_43_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_312_ _321_/CLK _312_/D VGND VGND VPWR VPWR _312_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_243_ _375_/CLK _243_/D VGND VGND VPWR VPWR _243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 a[25] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_4
X_174_ _319_/CLK _174_/D VGND VGND VPWR VPWR _174_/Q sky130_fd_sc_hd__dfxtp_1
Xinput29 a[35] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_93_2 dadda_fa_3_93_2/A dadda_fa_3_93_2/B dadda_fa_3_93_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_1/A dadda_fa_4_93_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_3_86_1 dadda_fa_3_86_1/A dadda_fa_3_86_1/B dadda_fa_3_86_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_0/CIN dadda_fa_4_86_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_63_0 dadda_fa_6_63_0/A dadda_fa_6_63_0/B dadda_fa_6_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_64_0/B dadda_fa_7_63_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_151_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_79_0 dadda_fa_3_79_0/A dadda_fa_3_79_0/B dadda_fa_3_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_0/B dadda_fa_4_79_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_ha_0_53_0 U$$113/X U$$246/X VGND VGND VPWR VPWR dadda_fa_1_54_8/B dadda_fa_2_53_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_42_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4301 U$$4438/A1 U$$4381/A2 U$$4440/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4302/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4312 U$$4312/A U$$4368/B VGND VGND VPWR VPWR U$$4312/X sky130_fd_sc_hd__xor2_1
XU$$4323 U$$4460/A1 U$$4349/A2 U$$4460/B1 U$$4349/B2 VGND VGND VPWR VPWR U$$4324/A
+ sky130_fd_sc_hd__a22o_1
XU$$4334 U$$4334/A U$$4360/B VGND VGND VPWR VPWR U$$4334/X sky130_fd_sc_hd__xor2_1
XU$$3600 U$$4420/B1 U$$3604/A2 U$$4287/A1 U$$3604/B2 VGND VGND VPWR VPWR U$$3601/A
+ sky130_fd_sc_hd__a22o_1
XU$$4345 U$$4345/A1 U$$4349/A2 U$$4482/B1 U$$4349/B2 VGND VGND VPWR VPWR U$$4346/A
+ sky130_fd_sc_hd__a22o_1
XU$$4356 U$$4356/A U$$4360/B VGND VGND VPWR VPWR U$$4356/X sky130_fd_sc_hd__xor2_1
XU$$3611 U$$3611/A U$$3615/B VGND VGND VPWR VPWR U$$3611/X sky130_fd_sc_hd__xor2_1
XU$$3622 U$$4307/A1 U$$3640/A2 U$$4307/B1 U$$3640/B2 VGND VGND VPWR VPWR U$$3623/A
+ sky130_fd_sc_hd__a22o_1
XU$$4367 U$$4504/A1 U$$4369/A2 U$$4367/B1 U$$4369/B2 VGND VGND VPWR VPWR U$$4368/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_115_1 U$$4360/X U$$4493/X input146/X VGND VGND VPWR VPWR dadda_fa_5_116_0/B
+ dadda_fa_5_115_1/B sky130_fd_sc_hd__fa_1
XU$$3633 U$$3633/A U$$3641/B VGND VGND VPWR VPWR U$$3633/X sky130_fd_sc_hd__xor2_1
XFILLER_19_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_867 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4378 U$$4378/A U$$4383/A VGND VGND VPWR VPWR U$$4378/X sky130_fd_sc_hd__xor2_1
XU$$4389 U$$4387/B U$$4384/A U$$4389/B1 U$$4384/Y VGND VGND VPWR VPWR U$$4389/X sky130_fd_sc_hd__a22o_4
XU$$3644 U$$4466/A1 U$$3644/A2 U$$4468/A1 U$$3644/B2 VGND VGND VPWR VPWR U$$3645/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3655 U$$3655/A U$$3659/B VGND VGND VPWR VPWR U$$3655/X sky130_fd_sc_hd__xor2_1
XU$$2910 U$$2910/A U$$2944/B VGND VGND VPWR VPWR U$$2910/X sky130_fd_sc_hd__xor2_1
XU$$3666 U$$4349/B1 U$$3682/A2 U$$4214/B1 U$$3682/B2 VGND VGND VPWR VPWR U$$3667/A
+ sky130_fd_sc_hd__a22o_1
XU$$2921 U$$3056/B1 U$$2937/A2 U$$2923/A1 U$$2937/B2 VGND VGND VPWR VPWR U$$2922/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_108_0 dadda_fa_4_108_0/A dadda_fa_4_108_0/B dadda_fa_4_108_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_109_0/A dadda_fa_5_108_1/A sky130_fd_sc_hd__fa_1
XU$$2932 U$$2932/A U$$2938/B VGND VGND VPWR VPWR U$$2932/X sky130_fd_sc_hd__xor2_1
XU$$3677 U$$3677/A U$$3698/A VGND VGND VPWR VPWR U$$3677/X sky130_fd_sc_hd__xor2_1
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2943 U$$612/B1 U$$2991/A2 U$$479/A1 U$$2991/B2 VGND VGND VPWR VPWR U$$2944/A sky130_fd_sc_hd__a22o_1
XU$$3688 U$$4508/B1 U$$3696/A2 U$$4375/A1 U$$3696/B2 VGND VGND VPWR VPWR U$$3689/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2954 U$$2954/A U$$3004/B VGND VGND VPWR VPWR U$$2954/X sky130_fd_sc_hd__xor2_1
XU$$3699 U$$3699/A VGND VGND VPWR VPWR U$$3699/Y sky130_fd_sc_hd__inv_1
XU$$2965 U$$3239/A1 U$$2979/A2 U$$3239/B1 U$$2979/B2 VGND VGND VPWR VPWR U$$2966/A
+ sky130_fd_sc_hd__a22o_1
XU$$2976 U$$2976/A U$$3014/A VGND VGND VPWR VPWR U$$2976/X sky130_fd_sc_hd__xor2_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2987 U$$4081/B1 U$$3005/A2 U$$3948/A1 U$$3005/B2 VGND VGND VPWR VPWR U$$2988/A
+ sky130_fd_sc_hd__a22o_1
XU$$2998 U$$2998/A U$$3004/B VGND VGND VPWR VPWR U$$2998/X sky130_fd_sc_hd__xor2_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4477_1886 VGND VGND VPWR VPWR U$$4477_1886/HI U$$4477/B sky130_fd_sc_hd__conb_1
Xdadda_fa_2_81_0 U$$4425/X input236/X dadda_fa_2_81_0/CIN VGND VGND VPWR VPWR dadda_fa_3_82_0/B
+ dadda_fa_3_81_2/B sky130_fd_sc_hd__fa_1
Xdadda_ha_1_51_8 U$$3301/X U$$3434/X VGND VGND VPWR VPWR dadda_fa_2_52_3/A dadda_fa_3_51_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_142_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$905 final_adder.U$$134/A final_adder.U$$843/X final_adder.U$$905/B1
+ VGND VGND VPWR VPWR final_adder.U$$905/X sky130_fd_sc_hd__a21o_1
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$927 final_adder.U$$156/A final_adder.U$$865/X final_adder.U$$927/B1
+ VGND VGND VPWR VPWR final_adder.U$$927/X sky130_fd_sc_hd__a21o_1
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$949 final_adder.U$$178/A final_adder.U$$887/X final_adder.U$$949/B1
+ VGND VGND VPWR VPWR final_adder.U$$949/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_6 U$$2501/X U$$2634/X U$$2767/X VGND VGND VPWR VPWR dadda_fa_2_51_2/B
+ dadda_fa_2_50_5/B sky130_fd_sc_hd__fa_1
XFILLER_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_2_0 U$$180/B input179/X dadda_ha_6_2_0/SUM VGND VGND VPWR VPWR _299_/D
+ _170_/D sky130_fd_sc_hd__fa_1
XFILLER_36_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_80_0 dadda_fa_7_80_0/A dadda_fa_7_80_0/B dadda_fa_7_80_0/CIN VGND VGND
+ VPWR VPWR _377_/D _248_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_96_0 dadda_fa_4_96_0/A dadda_fa_4_96_0/B dadda_fa_4_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_97_0/A dadda_fa_5_96_1/A sky130_fd_sc_hd__fa_1
XFILLER_146_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1105 U$$876/A1 VGND VGND VPWR VPWR U$$739/A1 sky130_fd_sc_hd__buf_4
Xfanout1116 U$$3751/A1 VGND VGND VPWR VPWR U$$4436/A1 sky130_fd_sc_hd__clkbuf_2
Xfanout1127 U$$2925/A1 VGND VGND VPWR VPWR U$$868/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1138 U$$8/B1 VGND VGND VPWR VPWR U$$10/A1 sky130_fd_sc_hd__buf_2
Xfanout1149 input75/X VGND VGND VPWR VPWR U$$4017/B1 sky130_fd_sc_hd__buf_6
XFILLER_87_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2206 U$$562/A1 U$$2248/A2 U$$562/B1 U$$2248/B2 VGND VGND VPWR VPWR U$$2207/A sky130_fd_sc_hd__a22o_1
XFILLER_170_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2217 U$$2217/A U$$2231/B VGND VGND VPWR VPWR U$$2217/X sky130_fd_sc_hd__xor2_1
XFILLER_74_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2228 U$$3322/B1 U$$2254/A2 U$$3189/A1 U$$2254/B2 VGND VGND VPWR VPWR U$$2229/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2239 U$$2239/A U$$2249/B VGND VGND VPWR VPWR U$$2239/X sky130_fd_sc_hd__xor2_1
XU$$1505 U$$1505/A U$$1507/A VGND VGND VPWR VPWR U$$1505/X sky130_fd_sc_hd__xor2_1
XU$$1516 U$$1516/A U$$1570/B VGND VGND VPWR VPWR U$$1516/X sky130_fd_sc_hd__xor2_1
XFILLER_103_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3294_1818 VGND VGND VPWR VPWR U$$3294_1818/HI U$$3294/A1 sky130_fd_sc_hd__conb_1
XU$$1527 U$$2758/B1 U$$1563/A2 U$$2625/A1 U$$1563/B2 VGND VGND VPWR VPWR U$$1528/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1538 U$$1538/A U$$1570/B VGND VGND VPWR VPWR U$$1538/X sky130_fd_sc_hd__xor2_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1549 U$$999/B1 U$$1567/A2 U$$866/A1 U$$1567/B2 VGND VGND VPWR VPWR U$$1550/A sky130_fd_sc_hd__a22o_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_226_ _356_/CLK _226_/D VGND VGND VPWR VPWR _226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_5 dadda_fa_2_60_5/A dadda_fa_2_60_5/B dadda_fa_2_60_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_2/A dadda_fa_4_60_0/A sky130_fd_sc_hd__fa_2
XFILLER_78_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1650 U$$4498/A1 VGND VGND VPWR VPWR U$$4361/A1 sky130_fd_sc_hd__buf_4
Xfanout1661 U$$4496/A1 VGND VGND VPWR VPWR U$$4359/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1672 input111/X VGND VGND VPWR VPWR U$$2711/B1 sky130_fd_sc_hd__buf_4
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4120 U$$4257/A1 U$$4158/A2 U$$4257/B1 U$$4158/B2 VGND VGND VPWR VPWR U$$4121/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_53_4 dadda_fa_2_53_4/A dadda_fa_2_53_4/B dadda_fa_2_53_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_1/CIN dadda_fa_3_53_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4131 U$$4131/A U$$4133/B VGND VGND VPWR VPWR U$$4131/X sky130_fd_sc_hd__xor2_1
Xfanout1683 U$$1328/B VGND VGND VPWR VPWR U$$1300/B sky130_fd_sc_hd__clkbuf_4
Xfanout1694 U$$3850/B1 VGND VGND VPWR VPWR U$$4400/A1 sky130_fd_sc_hd__buf_4
XU$$4142 U$$4416/A1 U$$4190/A2 U$$4416/B1 U$$4190/B2 VGND VGND VPWR VPWR U$$4143/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_46_3 dadda_fa_2_46_3/A dadda_fa_2_46_3/B dadda_fa_2_46_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_1/B dadda_fa_3_46_3/B sky130_fd_sc_hd__fa_1
XFILLER_65_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4153 U$$4153/A U$$4247/A VGND VGND VPWR VPWR U$$4153/X sky130_fd_sc_hd__xor2_1
XU$$4164 U$$4438/A1 U$$4174/A2 U$$4440/A1 U$$4174/B2 VGND VGND VPWR VPWR U$$4165/A
+ sky130_fd_sc_hd__a22o_1
XU$$4175 U$$4175/A U$$4175/B VGND VGND VPWR VPWR U$$4175/X sky130_fd_sc_hd__xor2_1
XFILLER_66_889 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3430 U$$3428/B U$$3425/A input46/X U$$3425/Y VGND VGND VPWR VPWR U$$3430/X sky130_fd_sc_hd__a22o_2
XU$$4186 U$$4460/A1 U$$4190/A2 U$$4460/B1 U$$4190/B2 VGND VGND VPWR VPWR U$$4187/A
+ sky130_fd_sc_hd__a22o_1
XU$$3441 U$$3713/B1 U$$3523/A2 U$$3580/A1 U$$3523/B2 VGND VGND VPWR VPWR U$$3442/A
+ sky130_fd_sc_hd__a22o_1
XU$$3452 U$$3452/A U$$3474/B VGND VGND VPWR VPWR U$$3452/X sky130_fd_sc_hd__xor2_1
XU$$4197 U$$4197/A U$$4215/B VGND VGND VPWR VPWR U$$4197/X sky130_fd_sc_hd__xor2_1
XU$$3463 U$$4420/B1 U$$3471/A2 U$$4287/A1 U$$3471/B2 VGND VGND VPWR VPWR U$$3464/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_39_2 U$$1947/X U$$2080/X U$$2213/X VGND VGND VPWR VPWR dadda_fa_3_40_1/A
+ dadda_fa_3_39_3/A sky130_fd_sc_hd__fa_1
XFILLER_129_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3474 U$$3474/A U$$3474/B VGND VGND VPWR VPWR U$$3474/X sky130_fd_sc_hd__xor2_1
XU$$2740 U$$2740/A VGND VGND VPWR VPWR U$$2740/Y sky130_fd_sc_hd__inv_1
XU$$3485 U$$4444/A1 U$$3557/A2 U$$4446/A1 U$$3557/B2 VGND VGND VPWR VPWR U$$3486/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_16_1 dadda_fa_5_16_1/A dadda_fa_5_16_1/B dadda_fa_5_16_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_17_0/B dadda_fa_7_16_0/A sky130_fd_sc_hd__fa_2
XU$$2751 U$$2751/A U$$2799/B VGND VGND VPWR VPWR U$$2751/X sky130_fd_sc_hd__xor2_1
XU$$3496 U$$3496/A U$$3506/B VGND VGND VPWR VPWR U$$3496/X sky130_fd_sc_hd__xor2_1
XU$$2762 U$$2897/B1 U$$2804/A2 U$$2762/B1 U$$2804/B2 VGND VGND VPWR VPWR U$$2763/A
+ sky130_fd_sc_hd__a22o_1
XU$$2773 U$$2773/A U$$2811/B VGND VGND VPWR VPWR U$$2773/X sky130_fd_sc_hd__xor2_1
XU$$2784 U$$866/A1 U$$2804/A2 U$$868/A1 U$$2804/B2 VGND VGND VPWR VPWR U$$2785/A sky130_fd_sc_hd__a22o_1
XU$$2795 U$$2795/A U$$2799/B VGND VGND VPWR VPWR U$$2795/X sky130_fd_sc_hd__xor2_1
XFILLER_167_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_42_4 U$$1687/X U$$1820/X VGND VGND VPWR VPWR dadda_fa_2_43_4/B dadda_fa_3_42_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_102_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput208 c[56] VGND VGND VPWR VPWR input208/X sky130_fd_sc_hd__clkbuf_4
Xinput219 c[66] VGND VGND VPWR VPWR input219/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$702 final_adder.U$$718/B final_adder.U$$702/B VGND VGND VPWR VPWR
+ final_adder.U$$782/A sky130_fd_sc_hd__and2_1
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$713 final_adder.U$$712/B final_adder.U$$609/X final_adder.U$$593/X
+ VGND VGND VPWR VPWR final_adder.U$$713/X sky130_fd_sc_hd__a21o_1
Xdadda_ha_4_12_2 U$$829/X U$$913/B VGND VGND VPWR VPWR dadda_fa_5_13_0/CIN dadda_ha_4_12_2/SUM
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$735 final_adder.U$$718/A final_adder.U$$381/X final_adder.U$$615/X
+ VGND VGND VPWR VPWR final_adder.U$$735/X sky130_fd_sc_hd__a21o_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$746 final_adder.U$$778/B final_adder.U$$746/B VGND VGND VPWR VPWR
+ final_adder.U$$746/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$757 final_adder.U$$756/B final_adder.U$$677/X final_adder.U$$645/X
+ VGND VGND VPWR VPWR final_adder.U$$757/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$768 final_adder.U$$800/B final_adder.U$$768/B VGND VGND VPWR VPWR
+ final_adder.U$$768/X sky130_fd_sc_hd__and2_1
XU$$607 U$$607/A U$$607/B VGND VGND VPWR VPWR U$$607/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$779 final_adder.U$$778/B final_adder.U$$699/X final_adder.U$$667/X
+ VGND VGND VPWR VPWR final_adder.U$$779/X sky130_fd_sc_hd__a21o_1
XFILLER_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$618 U$$892/A1 U$$636/A2 U$$894/A1 U$$636/B2 VGND VGND VPWR VPWR U$$619/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_41_2 U$$887/X U$$1020/X U$$1153/X VGND VGND VPWR VPWR dadda_fa_2_42_4/A
+ dadda_fa_2_41_5/CIN sky130_fd_sc_hd__fa_1
XU$$629 U$$629/A U$$631/B VGND VGND VPWR VPWR U$$629/X sky130_fd_sc_hd__xor2_1
XFILLER_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_11_0 U$$29/X U$$162/X U$$295/X VGND VGND VPWR VPWR dadda_fa_5_12_0/B dadda_fa_5_11_1/B
+ sky130_fd_sc_hd__fa_1
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_115_0 U$$3561/Y U$$3695/X U$$3828/X VGND VGND VPWR VPWR dadda_fa_4_116_2/B
+ dadda_fa_4_115_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_63_3 dadda_fa_3_63_3/A dadda_fa_3_63_3/B dadda_fa_3_63_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_1/B dadda_fa_4_63_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_56_2 dadda_fa_3_56_2/A dadda_fa_3_56_2/B dadda_fa_3_56_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_1/A dadda_fa_4_56_2/B sky130_fd_sc_hd__fa_1
XFILLER_47_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4387_1839 VGND VGND VPWR VPWR U$$4387_1839/HI U$$4387/A sky130_fd_sc_hd__conb_1
Xdadda_fa_3_49_1 dadda_fa_3_49_1/A dadda_fa_3_49_1/B dadda_fa_3_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_0/CIN dadda_fa_4_49_2/A sky130_fd_sc_hd__fa_1
XFILLER_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_26_0 dadda_fa_6_26_0/A dadda_fa_6_26_0/B dadda_fa_6_26_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_27_0/B dadda_fa_7_26_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_90_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2003 U$$2003/A U$$2031/B VGND VGND VPWR VPWR U$$2003/X sky130_fd_sc_hd__xor2_1
XFILLER_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2014 U$$918/A1 U$$2014/A2 U$$920/A1 U$$2014/B2 VGND VGND VPWR VPWR U$$2015/A sky130_fd_sc_hd__a22o_1
XU$$2025 U$$2025/A U$$2053/B VGND VGND VPWR VPWR U$$2025/X sky130_fd_sc_hd__xor2_1
XFILLER_16_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2036 U$$2310/A1 U$$2044/A2 U$$942/A1 U$$2044/B2 VGND VGND VPWR VPWR U$$2037/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1302 U$$1302/A U$$1328/B VGND VGND VPWR VPWR U$$1302/X sky130_fd_sc_hd__xor2_1
XU$$2047 U$$2047/A U$$2055/A VGND VGND VPWR VPWR U$$2047/X sky130_fd_sc_hd__xor2_1
XU$$1313 U$$80/A1 U$$1359/A2 U$$82/A1 U$$1359/B2 VGND VGND VPWR VPWR U$$1314/A sky130_fd_sc_hd__a22o_1
XU$$2058 U$$2192/A U$$2058/B VGND VGND VPWR VPWR U$$2058/X sky130_fd_sc_hd__and2_1
XU$$1324 U$$1324/A U$$1328/B VGND VGND VPWR VPWR U$$1324/X sky130_fd_sc_hd__xor2_1
XFILLER_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2069 U$$973/A1 U$$2107/A2 U$$973/B1 U$$2107/B2 VGND VGND VPWR VPWR U$$2070/A sky130_fd_sc_hd__a22o_1
XU$$1335 U$$924/A1 U$$1367/A2 U$$926/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1336/A sky130_fd_sc_hd__a22o_1
XU$$1346 U$$1346/A U$$1358/B VGND VGND VPWR VPWR U$$1346/X sky130_fd_sc_hd__xor2_1
XU$$1357 U$$946/A1 U$$1359/A2 U$$948/A1 U$$1359/B2 VGND VGND VPWR VPWR U$$1358/A sky130_fd_sc_hd__a22o_1
XU$$1368 U$$1368/A U$$1370/A VGND VGND VPWR VPWR U$$1368/X sky130_fd_sc_hd__xor2_1
XFILLER_15_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1379 U$$1379/A U$$1415/B VGND VGND VPWR VPWR U$$1379/X sky130_fd_sc_hd__xor2_1
XFILLER_31_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_209_ _338_/CLK _209_/D VGND VGND VPWR VPWR _209_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$1140 final_adder.U$$138/A final_adder.U$$847/X VGND VGND VPWR VPWR
+ output275/A sky130_fd_sc_hd__xor2_1
XFILLER_116_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1151 final_adder.U$$1151/A final_adder.U$$899/X VGND VGND VPWR VPWR
+ output287/A sky130_fd_sc_hd__xor2_4
XFILLER_129_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout909 U$$1218/B2 VGND VGND VPWR VPWR U$$1226/B2 sky130_fd_sc_hd__buf_6
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_51_1 dadda_fa_2_51_1/A dadda_fa_2_51_1/B dadda_fa_2_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_0/CIN dadda_fa_3_51_2/CIN sky130_fd_sc_hd__fa_1
Xfanout1480 U$$1721/B VGND VGND VPWR VPWR U$$1703/B sky130_fd_sc_hd__buf_6
Xfanout1491 input16/X VGND VGND VPWR VPWR U$$1618/B sky130_fd_sc_hd__buf_4
Xdadda_fa_2_44_0 U$$2356/X U$$2489/X U$$2622/X VGND VGND VPWR VPWR dadda_fa_3_45_0/B
+ dadda_fa_3_44_2/B sky130_fd_sc_hd__fa_1
XFILLER_94_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$20 _316_/Q _188_/Q VGND VGND VPWR VPWR final_adder.U$$235/A2 final_adder.U$$234/A
+ sky130_fd_sc_hd__ha_1
XFILLER_65_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$31 _327_/Q _199_/Q VGND VGND VPWR VPWR final_adder.U$$225/B1 final_adder.U$$224/B
+ sky130_fd_sc_hd__ha_1
XU$$3260 U$$3260/A U$$3284/B VGND VGND VPWR VPWR U$$3260/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$42 _338_/Q _210_/Q VGND VGND VPWR VPWR final_adder.U$$983/B1 final_adder.U$$212/A
+ sky130_fd_sc_hd__ha_1
XU$$3271 U$$3817/B1 U$$3285/A2 U$$4093/B1 U$$3285/B2 VGND VGND VPWR VPWR U$$3272/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$53 _349_/Q _221_/Q VGND VGND VPWR VPWR final_adder.U$$203/B1 final_adder.U$$202/B
+ sky130_fd_sc_hd__ha_1
XU$$3282 U$$3282/A U$$3284/B VGND VGND VPWR VPWR U$$3282/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$64 _360_/Q _232_/Q VGND VGND VPWR VPWR final_adder.U$$961/B1 final_adder.U$$190/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3293 U$$3291/B U$$3288/A input43/X U$$3288/Y VGND VGND VPWR VPWR U$$3293/X sky130_fd_sc_hd__a22o_4
Xfinal_adder.U$$75 _371_/Q _243_/Q VGND VGND VPWR VPWR final_adder.U$$181/B1 final_adder.U$$180/B
+ sky130_fd_sc_hd__ha_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2570 U$$2707/A1 U$$2574/A2 U$$2707/B1 U$$2574/B2 VGND VGND VPWR VPWR U$$2571/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$86 _382_/Q _254_/Q VGND VGND VPWR VPWR final_adder.U$$939/B1 final_adder.U$$168/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$97 _393_/Q _265_/Q VGND VGND VPWR VPWR final_adder.U$$159/B1 final_adder.U$$158/B
+ sky130_fd_sc_hd__ha_1
XFILLER_62_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2581 U$$2581/A U$$2591/B VGND VGND VPWR VPWR U$$2581/X sky130_fd_sc_hd__xor2_1
XU$$2592 U$$948/A1 U$$2598/A2 U$$950/A1 U$$2598/B2 VGND VGND VPWR VPWR U$$2593/A sky130_fd_sc_hd__a22o_1
XFILLER_55_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1880 U$$1880/A U$$1916/B VGND VGND VPWR VPWR U$$1880/X sky130_fd_sc_hd__xor2_1
XU$$1891 U$$4220/A1 U$$1891/A2 U$$4220/B1 U$$1891/B2 VGND VGND VPWR VPWR U$$1892/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_73_2 dadda_fa_4_73_2/A dadda_fa_4_73_2/B dadda_fa_4_73_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_74_0/CIN dadda_fa_5_73_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_150_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_89_2 U$$2579/X U$$2712/X U$$2845/X VGND VGND VPWR VPWR dadda_fa_2_90_4/B
+ dadda_fa_2_89_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_66_1 dadda_fa_4_66_1/A dadda_fa_4_66_1/B dadda_fa_4_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_67_0/B dadda_fa_5_66_1/B sky130_fd_sc_hd__fa_1
XFILLER_62_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_918 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_43_0 dadda_fa_7_43_0/A dadda_fa_7_43_0/B dadda_fa_7_43_0/CIN VGND VGND
+ VPWR VPWR _340_/D _211_/D sky130_fd_sc_hd__fa_2
XFILLER_103_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_59_0 dadda_fa_4_59_0/A dadda_fa_4_59_0/B dadda_fa_4_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_60_0/A dadda_fa_5_59_1/A sky130_fd_sc_hd__fa_1
XFILLER_131_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$510 final_adder.U$$518/B final_adder.U$$510/B VGND VGND VPWR VPWR
+ final_adder.U$$630/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$521 final_adder.U$$520/B final_adder.U$$405/X final_adder.U$$397/X
+ VGND VGND VPWR VPWR final_adder.U$$521/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$532 final_adder.U$$540/B final_adder.U$$532/B VGND VGND VPWR VPWR
+ final_adder.U$$652/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$543 final_adder.U$$542/B final_adder.U$$427/X final_adder.U$$419/X
+ VGND VGND VPWR VPWR final_adder.U$$543/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$554 final_adder.U$$562/B final_adder.U$$554/B VGND VGND VPWR VPWR
+ final_adder.U$$674/B sky130_fd_sc_hd__and2_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$565 final_adder.U$$564/B final_adder.U$$449/X final_adder.U$$441/X
+ VGND VGND VPWR VPWR final_adder.U$$565/X sky130_fd_sc_hd__a21o_1
XU$$404 U$$539/B1 U$$408/A2 U$$406/A1 U$$408/B2 VGND VGND VPWR VPWR U$$405/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$576 final_adder.U$$584/B final_adder.U$$576/B VGND VGND VPWR VPWR
+ final_adder.U$$696/B sky130_fd_sc_hd__and2_1
XU$$415 U$$413/Y U$$412/A U$$411/A U$$414/X U$$411/Y VGND VGND VPWR VPWR U$$415/X
+ sky130_fd_sc_hd__a32o_4
Xfinal_adder.U$$587 final_adder.U$$586/B final_adder.U$$471/X final_adder.U$$463/X
+ VGND VGND VPWR VPWR final_adder.U$$587/X sky130_fd_sc_hd__a21o_1
XFILLER_151_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$426 U$$426/A U$$448/B VGND VGND VPWR VPWR U$$426/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$598 final_adder.U$$606/B final_adder.U$$598/B VGND VGND VPWR VPWR
+ final_adder.U$$718/B sky130_fd_sc_hd__and2_1
XFILLER_71_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$437 U$$709/B1 U$$505/A2 U$$576/A1 U$$505/B2 VGND VGND VPWR VPWR U$$438/A sky130_fd_sc_hd__a22o_1
XFILLER_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$448 U$$448/A U$$448/B VGND VGND VPWR VPWR U$$448/X sky130_fd_sc_hd__xor2_1
XU$$459 U$$596/A1 U$$497/A2 U$$596/B1 U$$497/B2 VGND VGND VPWR VPWR U$$460/A sky130_fd_sc_hd__a22o_1
XFILLER_71_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_61_0 dadda_fa_3_61_0/A dadda_fa_3_61_0/B dadda_fa_3_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_0/B dadda_fa_4_61_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_77_0 U$$958/Y U$$1092/X U$$1225/X VGND VGND VPWR VPWR dadda_fa_1_78_8/CIN
+ dadda_fa_2_77_0/A sky130_fd_sc_hd__fa_2
XFILLER_0_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_976 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$960 input6/X VGND VGND VPWR VPWR U$$962/B sky130_fd_sc_hd__inv_1
Xdadda_ha_4_8_0 U$$23/X U$$156/X VGND VGND VPWR VPWR dadda_fa_5_9_1/B dadda_ha_4_8_0/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_90_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$971 U$$971/A1 U$$981/A2 U$$973/A1 U$$981/B2 VGND VGND VPWR VPWR U$$972/A sky130_fd_sc_hd__a22o_1
XU$$1110 U$$697/B1 U$$1174/A2 U$$975/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1111/A sky130_fd_sc_hd__a22o_1
XU$$1121 U$$1121/A U$$1195/B VGND VGND VPWR VPWR U$$1121/X sky130_fd_sc_hd__xor2_1
XU$$982 U$$982/A U$$982/B VGND VGND VPWR VPWR U$$982/X sky130_fd_sc_hd__xor2_1
XU$$1132 U$$995/A1 U$$1194/A2 U$$721/B1 U$$1194/B2 VGND VGND VPWR VPWR U$$1133/A sky130_fd_sc_hd__a22o_1
XU$$993 U$$993/A1 U$$997/A2 U$$995/A1 U$$997/B2 VGND VGND VPWR VPWR U$$994/A sky130_fd_sc_hd__a22o_1
XFILLER_44_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1143 U$$1143/A U$$1175/B VGND VGND VPWR VPWR U$$1143/X sky130_fd_sc_hd__xor2_1
XU$$1154 U$$58/A1 U$$1164/A2 U$$60/A1 U$$1164/B2 VGND VGND VPWR VPWR U$$1155/A sky130_fd_sc_hd__a22o_1
XU$$1165 U$$1165/A U$$1195/B VGND VGND VPWR VPWR U$$1165/X sky130_fd_sc_hd__xor2_1
XU$$1176 U$$80/A1 U$$1218/A2 U$$82/A1 U$$1218/B2 VGND VGND VPWR VPWR U$$1177/A sky130_fd_sc_hd__a22o_1
XU$$1187 U$$1187/A U$$1227/B VGND VGND VPWR VPWR U$$1187/X sky130_fd_sc_hd__xor2_1
XU$$1198 U$$924/A1 U$$1230/A2 U$$926/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1199/A sky130_fd_sc_hd__a22o_1
XFILLER_148_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_83_1 dadda_fa_5_83_1/A dadda_fa_5_83_1/B dadda_fa_5_83_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_84_0/B dadda_fa_7_83_0/A sky130_fd_sc_hd__fa_2
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_99_1 U$$2865/X U$$2998/X U$$3131/X VGND VGND VPWR VPWR dadda_fa_3_100_1/B
+ dadda_fa_3_99_3/A sky130_fd_sc_hd__fa_1
XFILLER_144_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_76_0 dadda_fa_5_76_0/A dadda_fa_5_76_0/B dadda_fa_5_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_77_0/A dadda_fa_6_76_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout706 U$$4190/B2 VGND VGND VPWR VPWR U$$4224/B2 sky130_fd_sc_hd__buf_4
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout717 U$$3978/X VGND VGND VPWR VPWR U$$4057/B2 sky130_fd_sc_hd__buf_6
Xfanout728 U$$3777/B2 VGND VGND VPWR VPWR U$$3739/B2 sky130_fd_sc_hd__buf_2
XFILLER_113_864 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_75_8 dadda_fa_1_75_8/A dadda_fa_1_75_8/B dadda_fa_1_75_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_76_3/A dadda_fa_3_75_0/A sky130_fd_sc_hd__fa_2
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 U$$3692/B2 VGND VGND VPWR VPWR U$$3696/B2 sky130_fd_sc_hd__buf_4
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_7 dadda_fa_1_68_7/A dadda_fa_1_68_7/B dadda_fa_1_68_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_69_2/CIN dadda_fa_2_68_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4116_1832 VGND VGND VPWR VPWR U$$4116_1832/HI U$$4116/A1 sky130_fd_sc_hd__conb_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3090 U$$3775/A1 U$$3108/A2 U$$3775/B1 U$$3108/B2 VGND VGND VPWR VPWR U$$3091/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_94_0 dadda_fa_1_94_0/A U$$2190/X U$$2323/X VGND VGND VPWR VPWR dadda_fa_2_95_5/B
+ dadda_fa_2_94_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_162_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$340 final_adder.U$$342/B final_adder.U$$340/B VGND VGND VPWR VPWR
+ final_adder.U$$466/B sky130_fd_sc_hd__and2_1
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$351 final_adder.U$$350/B final_adder.U$$225/X final_adder.U$$223/X
+ VGND VGND VPWR VPWR final_adder.U$$351/X sky130_fd_sc_hd__a21o_1
XFILLER_57_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$362 final_adder.U$$364/B final_adder.U$$362/B VGND VGND VPWR VPWR
+ final_adder.U$$488/B sky130_fd_sc_hd__and2_1
XFILLER_45_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$201 U$$884/B1 U$$219/A2 U$$64/B1 U$$219/B2 VGND VGND VPWR VPWR U$$202/A sky130_fd_sc_hd__a22o_1
XFILLER_73_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_106_0 dadda_fa_6_106_0/A dadda_fa_6_106_0/B dadda_fa_6_106_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_107_0/B dadda_fa_7_106_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$373 final_adder.U$$372/B final_adder.U$$247/X final_adder.U$$245/X
+ VGND VGND VPWR VPWR final_adder.U$$373/X sky130_fd_sc_hd__a21o_1
XU$$212 U$$212/A U$$214/B VGND VGND VPWR VPWR U$$212/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$384 final_adder.U$$388/B final_adder.U$$384/B VGND VGND VPWR VPWR
+ final_adder.U$$508/B sky130_fd_sc_hd__and2_1
XU$$223 U$$632/B1 U$$229/A2 U$$499/A1 U$$229/B2 VGND VGND VPWR VPWR U$$224/A sky130_fd_sc_hd__a22o_1
XFILLER_55_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$395 final_adder.U$$394/B final_adder.U$$273/X final_adder.U$$269/X
+ VGND VGND VPWR VPWR final_adder.U$$395/X sky130_fd_sc_hd__a21o_1
XU$$234 U$$234/A U$$273/A VGND VGND VPWR VPWR U$$234/X sky130_fd_sc_hd__xor2_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$245 U$$517/B1 U$$253/A2 U$$384/A1 U$$253/B2 VGND VGND VPWR VPWR U$$246/A sky130_fd_sc_hd__a22o_1
XU$$256 U$$256/A U$$260/B VGND VGND VPWR VPWR U$$256/X sky130_fd_sc_hd__xor2_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_26_3 dadda_fa_3_26_3/A dadda_fa_3_26_3/B dadda_fa_3_26_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_27_1/B dadda_fa_4_26_2/CIN sky130_fd_sc_hd__fa_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$267 U$$539/B1 U$$271/A2 U$$406/A1 U$$271/B2 VGND VGND VPWR VPWR U$$268/A sky130_fd_sc_hd__a22o_1
XFILLER_44_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$278 U$$276/Y U$$275/A U$$274/A U$$277/X U$$274/Y VGND VGND VPWR VPWR U$$278/X
+ sky130_fd_sc_hd__a32o_4
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$289 U$$289/A U$$313/B VGND VGND VPWR VPWR U$$289/X sky130_fd_sc_hd__xor2_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_93_0 dadda_fa_6_93_0/A dadda_fa_6_93_0/B dadda_fa_6_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_94_0/B dadda_fa_7_93_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_127_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$6 U$$6/A1 U$$8/A2 U$$8/A1 U$$8/B2 VGND VGND VPWR VPWR U$$7/A sky130_fd_sc_hd__a22o_1
XFILLER_126_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput309 output309/A VGND VGND VPWR VPWR o[31] sky130_fd_sc_hd__buf_2
XFILLER_153_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$790 U$$790/A U$$804/B VGND VGND VPWR VPWR U$$790/X sky130_fd_sc_hd__xor2_1
XFILLER_35_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3020_1814 VGND VGND VPWR VPWR U$$3020_1814/HI U$$3020/A1 sky130_fd_sc_hd__conb_1
XFILLER_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_110_0_1936 VGND VGND VPWR VPWR dadda_fa_3_110_0/A dadda_fa_3_110_0_1936/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_144_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_80_6 U$$3492/X U$$3625/X U$$3758/X VGND VGND VPWR VPWR dadda_fa_2_81_2/CIN
+ dadda_fa_2_80_5/B sky130_fd_sc_hd__fa_1
Xfanout503 U$$3245/A2 VGND VGND VPWR VPWR U$$3207/A2 sky130_fd_sc_hd__buf_4
Xfanout514 U$$3018/X VGND VGND VPWR VPWR U$$3112/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_73_5 U$$3877/X U$$4010/X U$$4143/X VGND VGND VPWR VPWR dadda_fa_2_74_2/A
+ dadda_fa_2_73_5/A sky130_fd_sc_hd__fa_1
Xfanout525 U$$2881/X VGND VGND VPWR VPWR U$$2989/A2 sky130_fd_sc_hd__buf_2
Xfanout536 U$$278/X VGND VGND VPWR VPWR U$$386/A2 sky130_fd_sc_hd__buf_6
XFILLER_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout547 U$$2607/X VGND VGND VPWR VPWR U$$2707/A2 sky130_fd_sc_hd__buf_4
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout558 fanout561/X VGND VGND VPWR VPWR U$$2548/A2 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_1_66_4 U$$4129/X U$$4262/X U$$4395/X VGND VGND VPWR VPWR dadda_fa_2_67_1/CIN
+ dadda_fa_2_66_4/CIN sky130_fd_sc_hd__fa_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout569 U$$2333/X VGND VGND VPWR VPWR U$$2463/A2 sky130_fd_sc_hd__buf_6
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_59_3 U$$2785/X U$$2918/X U$$3051/X VGND VGND VPWR VPWR dadda_fa_2_60_1/B
+ dadda_fa_2_59_4/B sky130_fd_sc_hd__fa_1
XFILLER_67_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_36_2 dadda_fa_4_36_2/A dadda_fa_4_36_2/B dadda_fa_4_36_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_37_0/CIN dadda_fa_5_36_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_29_1 dadda_fa_4_29_1/A dadda_fa_4_29_1/B dadda_fa_4_29_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_30_0/B dadda_fa_5_29_1/B sky130_fd_sc_hd__fa_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_190_ _321_/CLK _190_/D VGND VGND VPWR VPWR _190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_0_62_5 U$$2126/X U$$2259/X VGND VGND VPWR VPWR dadda_fa_1_63_7/A dadda_fa_2_62_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4505 U$$4505/A U$$4505/B VGND VGND VPWR VPWR U$$4505/X sky130_fd_sc_hd__xor2_1
XU$$4516 U$$4516/A1 U$$4388/X U$$545/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4517/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_0_61_3 U$$1326/X U$$1459/X U$$1592/X VGND VGND VPWR VPWR dadda_fa_1_62_6/CIN
+ dadda_fa_1_61_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$19 U$$19/A U$$9/B VGND VGND VPWR VPWR U$$19/X sky130_fd_sc_hd__xor2_1
XU$$3804 U$$3804/A U$$3816/B VGND VGND VPWR VPWR U$$3804/X sky130_fd_sc_hd__xor2_1
XU$$3815 U$$3815/A1 U$$3825/A2 U$$3817/A1 U$$3825/B2 VGND VGND VPWR VPWR U$$3816/A
+ sky130_fd_sc_hd__a22o_1
XU$$3826 U$$3826/A U$$3835/A VGND VGND VPWR VPWR U$$3826/X sky130_fd_sc_hd__xor2_1
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3837 input52/X VGND VGND VPWR VPWR U$$3839/B sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$170 final_adder.U$$170/A final_adder.U$$170/B VGND VGND VPWR VPWR
+ final_adder.U$$298/B sky130_fd_sc_hd__and2_1
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$181 final_adder.U$$180/B final_adder.U$$951/B1 final_adder.U$$181/B1
+ VGND VGND VPWR VPWR final_adder.U$$181/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_3_31_1 dadda_fa_3_31_1/A dadda_fa_3_31_1/B dadda_fa_3_31_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_32_0/CIN dadda_fa_4_31_2/A sky130_fd_sc_hd__fa_1
XU$$3848 U$$4257/B1 U$$3892/A2 U$$4259/B1 U$$3892/B2 VGND VGND VPWR VPWR U$$3849/A
+ sky130_fd_sc_hd__a22o_1
XU$$3859 U$$3859/A U$$3867/B VGND VGND VPWR VPWR U$$3859/X sky130_fd_sc_hd__xor2_1
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$192 final_adder.U$$192/A final_adder.U$$192/B VGND VGND VPWR VPWR
+ final_adder.U$$320/B sky130_fd_sc_hd__and2_1
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_24_0 U$$720/X U$$853/X U$$986/X VGND VGND VPWR VPWR dadda_fa_4_25_0/B
+ dadda_fa_4_24_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_388_ _388_/CLK _388_/D VGND VGND VPWR VPWR _388_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_90_5 dadda_fa_2_90_5/A dadda_fa_2_90_5/B dadda_fa_2_90_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_91_2/A dadda_fa_4_90_0/A sky130_fd_sc_hd__fa_2
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_83_4 dadda_fa_2_83_4/A dadda_fa_2_83_4/B dadda_fa_2_83_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_1/CIN dadda_fa_3_83_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_76_3 dadda_fa_2_76_3/A dadda_fa_2_76_3/B dadda_fa_2_76_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_1/B dadda_fa_3_76_3/B sky130_fd_sc_hd__fa_1
XFILLER_96_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_69_2 dadda_fa_2_69_2/A dadda_fa_2_69_2/B dadda_fa_2_69_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_1/A dadda_fa_3_69_3/A sky130_fd_sc_hd__fa_1
XFILLER_68_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_46_1 dadda_fa_5_46_1/A dadda_fa_5_46_1/B dadda_fa_5_46_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_47_0/B dadda_fa_7_46_0/A sky130_fd_sc_hd__fa_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_39_0 dadda_fa_5_39_0/A dadda_fa_5_39_0/B dadda_fa_5_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_40_0/A dadda_fa_6_39_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_64_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_120_1 dadda_fa_5_120_1/A dadda_fa_5_120_1/B dadda_ha_4_120_1/SUM VGND
+ VGND VPWR VPWR dadda_fa_6_121_0/B dadda_fa_7_120_0/A sky130_fd_sc_hd__fa_1
XFILLER_109_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_113_0 dadda_fa_5_113_0/A dadda_fa_5_113_0/B dadda_fa_5_113_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_114_0/A dadda_fa_6_113_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_137_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1309 input53/X VGND VGND VPWR VPWR fanout1309/X sky130_fd_sc_hd__buf_4
XFILLER_114_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_71_2 U$$2942/X U$$3075/X U$$3208/X VGND VGND VPWR VPWR dadda_fa_2_72_1/A
+ dadda_fa_2_71_4/A sky130_fd_sc_hd__fa_1
XFILLER_113_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_1 U$$2928/X U$$3061/X U$$3194/X VGND VGND VPWR VPWR dadda_fa_2_65_0/CIN
+ dadda_fa_2_64_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout388 U$$981/A2 VGND VGND VPWR VPWR U$$979/A2 sky130_fd_sc_hd__buf_4
Xfanout399 U$$826/X VGND VGND VPWR VPWR U$$952/A2 sky130_fd_sc_hd__buf_8
Xdadda_fa_4_41_0 dadda_fa_4_41_0/A dadda_fa_4_41_0/B dadda_fa_4_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_42_0/A dadda_fa_5_41_1/A sky130_fd_sc_hd__fa_1
XFILLER_28_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_57_0 U$$1185/X U$$1318/X U$$1451/X VGND VGND VPWR VPWR dadda_fa_2_58_0/B
+ dadda_fa_2_57_3/B sky130_fd_sc_hd__fa_1
XFILLER_46_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1709 U$$1709/A U$$1721/B VGND VGND VPWR VPWR U$$1709/X sky130_fd_sc_hd__xor2_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_311_ _321_/CLK _311_/D VGND VGND VPWR VPWR _311_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_242_ _247_/CLK _242_/D VGND VGND VPWR VPWR _242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_173_ _319_/CLK _173_/D VGND VGND VPWR VPWR _173_/Q sky130_fd_sc_hd__dfxtp_1
Xinput19 a[26] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_93_3 dadda_fa_3_93_3/A dadda_fa_3_93_3/B dadda_fa_3_93_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_1/B dadda_fa_4_93_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_124_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_86_2 dadda_fa_3_86_2/A dadda_fa_3_86_2/B dadda_fa_3_86_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_1/A dadda_fa_4_86_2/B sky130_fd_sc_hd__fa_1
XFILLER_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_79_1 dadda_fa_3_79_1/A dadda_fa_3_79_1/B dadda_fa_3_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_0/CIN dadda_fa_4_79_2/A sky130_fd_sc_hd__fa_1
XFILLER_96_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_56_0 dadda_fa_6_56_0/A dadda_fa_6_56_0/B dadda_fa_6_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_57_0/B dadda_fa_7_56_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_151_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4302 U$$4302/A U$$4384/A VGND VGND VPWR VPWR U$$4302/X sky130_fd_sc_hd__xor2_1
XFILLER_77_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4313 U$$4450/A1 U$$4373/A2 U$$4315/A1 U$$4373/B2 VGND VGND VPWR VPWR U$$4314/A
+ sky130_fd_sc_hd__a22o_1
XU$$4324 U$$4324/A U$$4350/B VGND VGND VPWR VPWR U$$4324/X sky130_fd_sc_hd__xor2_1
XU$$4335 U$$4472/A1 U$$4349/A2 U$$4474/A1 U$$4349/B2 VGND VGND VPWR VPWR U$$4336/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3601 U$$3601/A U$$3601/B VGND VGND VPWR VPWR U$$3601/X sky130_fd_sc_hd__xor2_1
XU$$4346 U$$4346/A U$$4350/B VGND VGND VPWR VPWR U$$4346/X sky130_fd_sc_hd__xor2_1
XU$$4357 U$$4492/B1 U$$4359/A2 U$$4359/A1 U$$4359/B2 VGND VGND VPWR VPWR U$$4358/A
+ sky130_fd_sc_hd__a22o_1
XU$$3612 U$$4434/A1 U$$3656/A2 U$$3751/A1 U$$3656/B2 VGND VGND VPWR VPWR U$$3613/A
+ sky130_fd_sc_hd__a22o_1
XU$$3623 U$$3623/A U$$3641/B VGND VGND VPWR VPWR U$$3623/X sky130_fd_sc_hd__xor2_1
XU$$4368 U$$4368/A U$$4368/B VGND VGND VPWR VPWR U$$4368/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_115_2 dadda_fa_4_115_2/A dadda_fa_4_115_2/B dadda_fa_4_115_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_116_0/CIN dadda_fa_5_115_1/CIN sky130_fd_sc_hd__fa_1
XU$$3634 U$$4043/B1 U$$3640/A2 U$$3908/B1 U$$3640/B2 VGND VGND VPWR VPWR U$$3635/A
+ sky130_fd_sc_hd__a22o_1
XU$$4379 U$$4516/A1 U$$4381/A2 U$$545/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4380/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3645 U$$3645/A U$$3699/A VGND VGND VPWR VPWR U$$3645/X sky130_fd_sc_hd__xor2_1
XU$$2900 U$$2900/A U$$2944/B VGND VGND VPWR VPWR U$$2900/X sky130_fd_sc_hd__xor2_1
XFILLER_80_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3656 U$$4478/A1 U$$3656/A2 U$$4478/B1 U$$3656/B2 VGND VGND VPWR VPWR U$$3657/A
+ sky130_fd_sc_hd__a22o_1
XU$$2911 U$$3048/A1 U$$2991/A2 U$$3048/B1 U$$2991/B2 VGND VGND VPWR VPWR U$$2912/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2922 U$$2922/A U$$2938/B VGND VGND VPWR VPWR U$$2922/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_108_1 dadda_fa_4_108_1/A dadda_fa_4_108_1/B dadda_fa_4_108_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_109_0/B dadda_fa_5_108_1/B sky130_fd_sc_hd__fa_1
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3667 U$$3667/A U$$3681/B VGND VGND VPWR VPWR U$$3667/X sky130_fd_sc_hd__xor2_1
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2933 U$$4027/B1 U$$2937/A2 U$$4442/A1 U$$2937/B2 VGND VGND VPWR VPWR U$$2934/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3678 U$$3815/A1 U$$3682/A2 U$$3817/A1 U$$3682/B2 VGND VGND VPWR VPWR U$$3679/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2944 U$$2944/A U$$2944/B VGND VGND VPWR VPWR U$$2944/X sky130_fd_sc_hd__xor2_1
XU$$3689 U$$3689/A U$$3695/B VGND VGND VPWR VPWR U$$3689/X sky130_fd_sc_hd__xor2_1
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2955 U$$4462/A1 U$$3011/A2 U$$3916/A1 U$$3011/B2 VGND VGND VPWR VPWR U$$2956/A
+ sky130_fd_sc_hd__a22o_1
XU$$2966 U$$2966/A U$$2974/B VGND VGND VPWR VPWR U$$2966/X sky130_fd_sc_hd__xor2_1
XU$$2977 U$$922/A1 U$$2977/A2 U$$922/B1 U$$2977/B2 VGND VGND VPWR VPWR U$$2978/A sky130_fd_sc_hd__a22o_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2988 U$$2988/A U$$3004/B VGND VGND VPWR VPWR U$$2988/X sky130_fd_sc_hd__xor2_1
XU$$2999 U$$3684/A1 U$$3011/A2 U$$3684/B1 U$$3011/B2 VGND VGND VPWR VPWR U$$3000/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_81_1 dadda_fa_2_81_1/A dadda_fa_2_81_1/B dadda_fa_2_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_0/CIN dadda_fa_3_81_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_138_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_74_0 dadda_fa_2_74_0/A dadda_fa_2_74_0/B dadda_fa_2_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_0/B dadda_fa_3_74_2/B sky130_fd_sc_hd__fa_1
XFILLER_69_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$917 final_adder.U$$146/A final_adder.U$$855/X final_adder.U$$917/B1
+ VGND VGND VPWR VPWR final_adder.U$$917/X sky130_fd_sc_hd__a21o_1
XFILLER_29_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$939 final_adder.U$$168/A final_adder.U$$877/X final_adder.U$$939/B1
+ VGND VGND VPWR VPWR final_adder.U$$939/X sky130_fd_sc_hd__a21o_1
XFILLER_83_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_50_7 U$$2900/X U$$3033/X U$$3166/X VGND VGND VPWR VPWR dadda_fa_2_51_2/CIN
+ dadda_fa_2_50_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_96_1 dadda_fa_4_96_1/A dadda_fa_4_96_1/B dadda_fa_4_96_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_97_0/B dadda_fa_5_96_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_7_73_0 dadda_fa_7_73_0/A dadda_fa_7_73_0/B dadda_fa_7_73_0/CIN VGND VGND
+ VPWR VPWR _370_/D _241_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_89_0 dadda_fa_4_89_0/A dadda_fa_4_89_0/B dadda_fa_4_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_90_0/A dadda_fa_5_89_1/A sky130_fd_sc_hd__fa_1
XFILLER_152_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1106 input80/X VGND VGND VPWR VPWR U$$876/A1 sky130_fd_sc_hd__buf_6
Xfanout1117 input79/X VGND VGND VPWR VPWR U$$3751/A1 sky130_fd_sc_hd__buf_4
Xfanout1128 U$$3884/A1 VGND VGND VPWR VPWR U$$2925/A1 sky130_fd_sc_hd__buf_4
Xfanout1139 U$$3435/A1 VGND VGND VPWR VPWR U$$8/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2207 U$$2207/A U$$2253/B VGND VGND VPWR VPWR U$$2207/X sky130_fd_sc_hd__xor2_1
XU$$2218 U$$983/B1 U$$2254/A2 U$$850/A1 U$$2254/B2 VGND VGND VPWR VPWR U$$2219/A sky130_fd_sc_hd__a22o_1
XU$$2229 U$$2229/A U$$2231/B VGND VGND VPWR VPWR U$$2229/X sky130_fd_sc_hd__xor2_1
XFILLER_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1506 U$$1507/A VGND VGND VPWR VPWR U$$1506/Y sky130_fd_sc_hd__inv_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1517 U$$3296/B1 U$$1567/A2 U$$3298/B1 U$$1567/B2 VGND VGND VPWR VPWR U$$1518/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1528 U$$1528/A U$$1564/B VGND VGND VPWR VPWR U$$1528/X sky130_fd_sc_hd__xor2_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1539 U$$32/A1 U$$1575/A2 U$$32/B1 U$$1575/B2 VGND VGND VPWR VPWR U$$1540/A sky130_fd_sc_hd__a22o_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_225_ _356_/CLK _225_/D VGND VGND VPWR VPWR _225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_91_0 dadda_fa_3_91_0/A dadda_fa_3_91_0/B dadda_fa_3_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_0/B dadda_fa_4_91_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_109_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1640 input114/X VGND VGND VPWR VPWR U$$253/A1 sky130_fd_sc_hd__buf_6
Xfanout1651 U$$4498/A1 VGND VGND VPWR VPWR U$$3948/B1 sky130_fd_sc_hd__buf_4
XFILLER_78_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4110 U$$4110/A VGND VGND VPWR VPWR U$$4110/Y sky130_fd_sc_hd__inv_1
Xfanout1662 U$$2578/A1 VGND VGND VPWR VPWR U$$4496/A1 sky130_fd_sc_hd__buf_2
XFILLER_93_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_120_0 dadda_fa_4_120_0/A U$$3971/X U$$4104/X VGND VGND VPWR VPWR dadda_fa_5_121_1/A
+ dadda_fa_5_120_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_2_53_5 dadda_fa_2_53_5/A dadda_fa_2_53_5/B dadda_fa_2_53_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_2/A dadda_fa_4_53_0/A sky130_fd_sc_hd__fa_1
XU$$4121 U$$4121/A U$$4133/B VGND VGND VPWR VPWR U$$4121/X sky130_fd_sc_hd__xor2_1
Xfanout1673 U$$2711/A1 VGND VGND VPWR VPWR U$$2574/A1 sky130_fd_sc_hd__buf_4
Xfanout1684 U$$1360/B VGND VGND VPWR VPWR U$$1328/B sky130_fd_sc_hd__buf_6
XU$$4132 U$$4132/A1 U$$4158/A2 U$$4132/B1 U$$4158/B2 VGND VGND VPWR VPWR U$$4133/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1695 input109/X VGND VGND VPWR VPWR U$$3850/B1 sky130_fd_sc_hd__buf_4
XFILLER_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4143 U$$4143/A U$$4191/B VGND VGND VPWR VPWR U$$4143/X sky130_fd_sc_hd__xor2_1
XU$$4154 U$$4291/A1 U$$4174/A2 U$$4291/B1 U$$4174/B2 VGND VGND VPWR VPWR U$$4155/A
+ sky130_fd_sc_hd__a22o_1
XU$$4165 U$$4165/A U$$4175/B VGND VGND VPWR VPWR U$$4165/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_46_4 dadda_fa_2_46_4/A dadda_fa_2_46_4/B dadda_fa_2_46_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_1/CIN dadda_fa_3_46_3/CIN sky130_fd_sc_hd__fa_1
XU$$3420 U$$3966/B1 U$$3422/A2 U$$3833/A1 U$$3422/B2 VGND VGND VPWR VPWR U$$3421/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3431 U$$3431/A1 U$$3471/A2 U$$3979/B1 U$$3471/B2 VGND VGND VPWR VPWR U$$3432/A
+ sky130_fd_sc_hd__a22o_1
XU$$4176 U$$4176/A1 U$$4244/A2 U$$4176/B1 U$$4244/B2 VGND VGND VPWR VPWR U$$4177/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4187 U$$4187/A U$$4191/B VGND VGND VPWR VPWR U$$4187/X sky130_fd_sc_hd__xor2_1
XU$$3442 U$$3442/A U$$3482/B VGND VGND VPWR VPWR U$$3442/X sky130_fd_sc_hd__xor2_1
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3453 U$$3999/B1 U$$3471/A2 U$$4001/B1 U$$3471/B2 VGND VGND VPWR VPWR U$$3454/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4198 U$$4472/A1 U$$4224/A2 U$$4198/B1 U$$4224/B2 VGND VGND VPWR VPWR U$$4199/A
+ sky130_fd_sc_hd__a22o_1
XU$$3464 U$$3464/A U$$3468/B VGND VGND VPWR VPWR U$$3464/X sky130_fd_sc_hd__xor2_1
XFILLER_81_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_39_3 U$$2346/X U$$2479/X U$$2612/X VGND VGND VPWR VPWR dadda_fa_3_40_1/B
+ dadda_fa_3_39_3/B sky130_fd_sc_hd__fa_1
XU$$2730 U$$2730/A U$$2738/B VGND VGND VPWR VPWR U$$2730/X sky130_fd_sc_hd__xor2_1
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3475 U$$3610/B1 U$$3523/A2 U$$874/A1 U$$3523/B2 VGND VGND VPWR VPWR U$$3476/A
+ sky130_fd_sc_hd__a22o_1
XU$$2741 input35/X VGND VGND VPWR VPWR U$$2743/B sky130_fd_sc_hd__inv_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3486 U$$3486/A U$$3558/B VGND VGND VPWR VPWR U$$3486/X sky130_fd_sc_hd__xor2_1
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2752 U$$2887/B1 U$$2798/A2 U$$2754/A1 U$$2798/B2 VGND VGND VPWR VPWR U$$2753/A
+ sky130_fd_sc_hd__a22o_1
XU$$3497 U$$4043/B1 U$$3505/A2 U$$3499/A1 U$$3505/B2 VGND VGND VPWR VPWR U$$3498/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2763 U$$2763/A U$$2805/B VGND VGND VPWR VPWR U$$2763/X sky130_fd_sc_hd__xor2_1
XU$$2774 U$$32/B1 U$$2812/A2 U$$447/A1 U$$2812/B2 VGND VGND VPWR VPWR U$$2775/A sky130_fd_sc_hd__a22o_1
XU$$2785 U$$2785/A U$$2805/B VGND VGND VPWR VPWR U$$2785/X sky130_fd_sc_hd__xor2_1
XU$$2796 U$$4027/B1 U$$2840/A2 U$$4442/A1 U$$2840/B2 VGND VGND VPWR VPWR U$$2797/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput209 c[57] VGND VGND VPWR VPWR input209/X sky130_fd_sc_hd__buf_2
XFILLER_130_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$703 final_adder.U$$702/B final_adder.U$$599/X final_adder.U$$583/X
+ VGND VGND VPWR VPWR final_adder.U$$703/X sky130_fd_sc_hd__a21o_1
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$714 final_adder.U$$714/A final_adder.U$$714/B VGND VGND VPWR VPWR
+ final_adder.U$$794/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$725 final_adder.U$$708/A final_adder.U$$621/X final_adder.U$$605/X
+ VGND VGND VPWR VPWR final_adder.U$$725/X sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$747 final_adder.U$$746/B final_adder.U$$667/X final_adder.U$$635/X
+ VGND VGND VPWR VPWR final_adder.U$$747/X sky130_fd_sc_hd__a21o_1
XFILLER_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$758 final_adder.U$$790/B final_adder.U$$758/B VGND VGND VPWR VPWR
+ final_adder.U$$758/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$769 final_adder.U$$768/B final_adder.U$$689/X final_adder.U$$657/X
+ VGND VGND VPWR VPWR final_adder.U$$769/X sky130_fd_sc_hd__a21o_1
XFILLER_112_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$608 U$$882/A1 U$$642/A2 U$$882/B1 U$$642/B2 VGND VGND VPWR VPWR U$$609/A sky130_fd_sc_hd__a22o_1
XU$$619 U$$619/A U$$637/B VGND VGND VPWR VPWR U$$619/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_108_0 U$$3282/X U$$3415/X U$$3548/X VGND VGND VPWR VPWR dadda_fa_4_109_0/B
+ dadda_fa_4_108_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_56_3 dadda_fa_3_56_3/A dadda_fa_3_56_3/B dadda_fa_3_56_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_1/B dadda_fa_4_56_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_49_2 dadda_fa_3_49_2/A dadda_fa_3_49_2/B dadda_fa_3_49_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_1/A dadda_fa_4_49_2/B sky130_fd_sc_hd__fa_1
XFILLER_114_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2004 U$$3509/B1 U$$2046/A2 U$$3376/A1 U$$2046/B2 VGND VGND VPWR VPWR U$$2005/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2015 U$$2015/A U$$2015/B VGND VGND VPWR VPWR U$$2015/X sky130_fd_sc_hd__xor2_1
XU$$2026 U$$2574/A1 U$$2046/A2 U$$2576/A1 U$$2046/B2 VGND VGND VPWR VPWR U$$2027/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_19_0 dadda_fa_6_19_0/A dadda_fa_6_19_0/B dadda_fa_6_19_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_20_0/B dadda_fa_7_19_0/CIN sky130_fd_sc_hd__fa_1
XU$$2037 U$$2037/A U$$2043/B VGND VGND VPWR VPWR U$$2037/X sky130_fd_sc_hd__xor2_1
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2048 U$$4375/B1 U$$2052/A2 U$$4240/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2049/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1303 U$$481/A1 U$$1311/A2 U$$72/A1 U$$1311/B2 VGND VGND VPWR VPWR U$$1304/A sky130_fd_sc_hd__a22o_1
XU$$2059 U$$2057/Y input24/X U$$2055/A U$$2058/X U$$2055/Y VGND VGND VPWR VPWR U$$2059/X
+ sky130_fd_sc_hd__a32o_4
XU$$1314 U$$1314/A U$$1358/B VGND VGND VPWR VPWR U$$1314/X sky130_fd_sc_hd__xor2_1
XU$$1325 U$$92/A1 U$$1367/A2 U$$94/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1326/A sky130_fd_sc_hd__a22o_1
XU$$1336 U$$1336/A U$$1364/B VGND VGND VPWR VPWR U$$1336/X sky130_fd_sc_hd__xor2_1
XFILLER_128_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1347 U$$386/B1 U$$1359/A2 U$$253/A1 U$$1359/B2 VGND VGND VPWR VPWR U$$1348/A sky130_fd_sc_hd__a22o_1
XU$$1358 U$$1358/A U$$1358/B VGND VGND VPWR VPWR U$$1358/X sky130_fd_sc_hd__xor2_1
XU$$1369 U$$1370/A VGND VGND VPWR VPWR U$$1369/Y sky130_fd_sc_hd__inv_1
XFILLER_168_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_208_ _344_/CLK _208_/D VGND VGND VPWR VPWR _208_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$1130 final_adder.U$$148/A final_adder.U$$857/X VGND VGND VPWR VPWR
+ output264/A sky130_fd_sc_hd__xor2_1
XFILLER_157_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1141 final_adder.U$$138/B final_adder.U$$909/X VGND VGND VPWR VPWR
+ output276/A sky130_fd_sc_hd__xor2_1
XFILLER_8_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1470 U$$1854/B VGND VGND VPWR VPWR U$$1836/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_51_2 dadda_fa_2_51_2/A dadda_fa_2_51_2/B dadda_fa_2_51_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_1/A dadda_fa_3_51_3/A sky130_fd_sc_hd__fa_1
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1481 input18/X VGND VGND VPWR VPWR U$$1721/B sky130_fd_sc_hd__buf_6
XFILLER_65_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1492 U$$1630/B VGND VGND VPWR VPWR U$$1644/A sky130_fd_sc_hd__buf_6
Xdadda_fa_2_44_1 U$$2755/X U$$2888/X U$$3021/X VGND VGND VPWR VPWR dadda_fa_3_45_0/CIN
+ dadda_fa_3_44_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_94_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$10 _306_/Q _178_/Q VGND VGND VPWR VPWR final_adder.U$$245/A2 final_adder.U$$244/A
+ sky130_fd_sc_hd__ha_1
XFILLER_26_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$21 _317_/Q _189_/Q VGND VGND VPWR VPWR final_adder.U$$235/B1 final_adder.U$$234/B
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3250 U$$3250/A U$$3287/A VGND VGND VPWR VPWR U$$3250/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_21_0 dadda_fa_5_21_0/A dadda_fa_5_21_0/B dadda_fa_5_21_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_22_0/A dadda_fa_6_21_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$32 _328_/Q _200_/Q VGND VGND VPWR VPWR final_adder.U$$993/B1 final_adder.U$$222/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_2_37_0 U$$746/X U$$879/X U$$1012/X VGND VGND VPWR VPWR dadda_fa_3_38_0/B
+ dadda_fa_3_37_2/B sky130_fd_sc_hd__fa_1
XU$$3261 U$$4081/B1 U$$3283/A2 U$$3948/A1 U$$3283/B2 VGND VGND VPWR VPWR U$$3262/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$43 _339_/Q _211_/Q VGND VGND VPWR VPWR final_adder.U$$213/B1 final_adder.U$$212/B
+ sky130_fd_sc_hd__ha_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3272 U$$3272/A U$$3286/B VGND VGND VPWR VPWR U$$3272/X sky130_fd_sc_hd__xor2_1
XFILLER_80_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_94_0_1930 VGND VGND VPWR VPWR dadda_fa_1_94_0/A dadda_fa_1_94_0_1930/LO
+ sky130_fd_sc_hd__conb_1
Xfinal_adder.U$$54 _350_/Q _222_/Q VGND VGND VPWR VPWR final_adder.U$$971/B1 final_adder.U$$200/A
+ sky130_fd_sc_hd__ha_1
XU$$3283 U$$3418/B1 U$$3283/A2 U$$3285/A1 U$$3283/B2 VGND VGND VPWR VPWR U$$3284/A
+ sky130_fd_sc_hd__a22o_1
XU$$3294 U$$3294/A1 U$$3338/A2 U$$4392/A1 U$$3338/B2 VGND VGND VPWR VPWR U$$3295/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$65 _361_/Q _233_/Q VGND VGND VPWR VPWR final_adder.U$$191/B1 final_adder.U$$190/B
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$76 _372_/Q _244_/Q VGND VGND VPWR VPWR final_adder.U$$949/B1 final_adder.U$$178/A
+ sky130_fd_sc_hd__ha_1
XU$$2560 U$$3243/B1 U$$2574/A2 U$$3110/A1 U$$2574/B2 VGND VGND VPWR VPWR U$$2561/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$87 _383_/Q _255_/Q VGND VGND VPWR VPWR final_adder.U$$169/B1 final_adder.U$$168/B
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$98 _394_/Q _266_/Q VGND VGND VPWR VPWR final_adder.U$$927/B1 final_adder.U$$156/A
+ sky130_fd_sc_hd__ha_1
XU$$2571 U$$2571/A U$$2575/B VGND VGND VPWR VPWR U$$2571/X sky130_fd_sc_hd__xor2_1
XU$$2582 U$$4363/A1 U$$2598/A2 U$$4365/A1 U$$2598/B2 VGND VGND VPWR VPWR U$$2583/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2593 U$$2593/A U$$2602/A VGND VGND VPWR VPWR U$$2593/X sky130_fd_sc_hd__xor2_1
XU$$1870 U$$1870/A U$$1874/B VGND VGND VPWR VPWR U$$1870/X sky130_fd_sc_hd__xor2_1
XFILLER_142_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1881 U$$920/B1 U$$1881/A2 U$$787/A1 U$$1881/B2 VGND VGND VPWR VPWR U$$1882/A sky130_fd_sc_hd__a22o_1
XU$$1892 U$$1892/A U$$1916/B VGND VGND VPWR VPWR U$$1892/X sky130_fd_sc_hd__xor2_1
XFILLER_166_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_89_3 U$$2978/X U$$3111/X U$$3244/X VGND VGND VPWR VPWR dadda_fa_2_90_4/CIN
+ dadda_fa_3_89_0/A sky130_fd_sc_hd__fa_1
XFILLER_103_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_66_2 dadda_fa_4_66_2/A dadda_fa_4_66_2/B dadda_fa_4_66_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_67_0/CIN dadda_fa_5_66_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_59_1 dadda_fa_4_59_1/A dadda_fa_4_59_1/B dadda_fa_4_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_60_0/B dadda_fa_5_59_1/B sky130_fd_sc_hd__fa_1
XFILLER_130_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$500 final_adder.U$$500/A final_adder.U$$500/B VGND VGND VPWR VPWR
+ final_adder.U$$616/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$511 final_adder.U$$510/B final_adder.U$$395/X final_adder.U$$387/X
+ VGND VGND VPWR VPWR final_adder.U$$511/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_0_68_0_1918 VGND VGND VPWR VPWR dadda_fa_0_68_0/A dadda_fa_0_68_0_1918/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_85_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_36_0 dadda_fa_7_36_0/A dadda_fa_7_36_0/B dadda_fa_7_36_0/CIN VGND VGND
+ VPWR VPWR _333_/D _204_/D sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$522 final_adder.U$$530/B final_adder.U$$522/B VGND VGND VPWR VPWR
+ final_adder.U$$642/B sky130_fd_sc_hd__and2_1
XFILLER_28_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$533 final_adder.U$$532/B final_adder.U$$417/X final_adder.U$$409/X
+ VGND VGND VPWR VPWR final_adder.U$$533/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$544 final_adder.U$$552/B final_adder.U$$544/B VGND VGND VPWR VPWR
+ final_adder.U$$664/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$555 final_adder.U$$554/B final_adder.U$$439/X final_adder.U$$431/X
+ VGND VGND VPWR VPWR final_adder.U$$555/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$566 final_adder.U$$574/B final_adder.U$$566/B VGND VGND VPWR VPWR
+ final_adder.U$$686/B sky130_fd_sc_hd__and2_1
XU$$405 U$$405/A U$$411/A VGND VGND VPWR VPWR U$$405/X sky130_fd_sc_hd__xor2_1
XFILLER_56_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$577 final_adder.U$$576/B final_adder.U$$461/X final_adder.U$$453/X
+ VGND VGND VPWR VPWR final_adder.U$$577/X sky130_fd_sc_hd__a21o_1
XU$$416 U$$414/B U$$411/A U$$412/A U$$411/Y VGND VGND VPWR VPWR U$$416/X sky130_fd_sc_hd__a22o_4
Xfinal_adder.U$$588 final_adder.U$$596/B final_adder.U$$588/B VGND VGND VPWR VPWR
+ final_adder.U$$708/B sky130_fd_sc_hd__and2_1
XU$$427 U$$16/A1 U$$447/A2 U$$566/A1 U$$447/B2 VGND VGND VPWR VPWR U$$428/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$599 final_adder.U$$598/B final_adder.U$$483/X final_adder.U$$475/X
+ VGND VGND VPWR VPWR final_adder.U$$599/X sky130_fd_sc_hd__a21o_1
XFILLER_45_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$438 U$$438/A U$$506/B VGND VGND VPWR VPWR U$$438/X sky130_fd_sc_hd__xor2_1
XFILLER_151_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$449 U$$38/A1 U$$505/A2 U$$40/A1 U$$505/B2 VGND VGND VPWR VPWR U$$450/A sky130_fd_sc_hd__a22o_1
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4393_1844 VGND VGND VPWR VPWR U$$4393_1844/HI U$$4393/B sky130_fd_sc_hd__conb_1
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_61_1 dadda_fa_3_61_1/A dadda_fa_3_61_1/B dadda_fa_3_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_0/CIN dadda_fa_4_61_2/A sky130_fd_sc_hd__fa_1
XFILLER_79_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_54_0 dadda_fa_3_54_0/A dadda_fa_3_54_0/B dadda_fa_3_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_0/B dadda_fa_4_54_1/CIN sky130_fd_sc_hd__fa_1
Xclkbuf_2_3__f_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _370_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$950 U$$950/A1 U$$956/A2 U$$952/A1 U$$956/B2 VGND VGND VPWR VPWR U$$951/A sky130_fd_sc_hd__a22o_1
XU$$1100 U$$1098/Y input8/X U$$962/A U$$1099/X U$$1096/Y VGND VGND VPWR VPWR U$$1100/X
+ sky130_fd_sc_hd__a32o_1
XU$$961 U$$962/A VGND VGND VPWR VPWR U$$961/Y sky130_fd_sc_hd__inv_1
XFILLER_91_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$972 U$$972/A U$$982/B VGND VGND VPWR VPWR U$$972/X sky130_fd_sc_hd__xor2_1
XU$$1111 U$$1111/A U$$1175/B VGND VGND VPWR VPWR U$$1111/X sky130_fd_sc_hd__xor2_1
XU$$1122 U$$983/B1 U$$1164/A2 U$$850/A1 U$$1164/B2 VGND VGND VPWR VPWR U$$1123/A sky130_fd_sc_hd__a22o_1
XU$$983 U$$983/A1 U$$997/A2 U$$983/B1 U$$997/B2 VGND VGND VPWR VPWR U$$984/A sky130_fd_sc_hd__a22o_1
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$994 U$$994/A U$$998/B VGND VGND VPWR VPWR U$$994/X sky130_fd_sc_hd__xor2_1
XU$$1133 U$$1133/A U$$1195/B VGND VGND VPWR VPWR U$$1133/X sky130_fd_sc_hd__xor2_1
XFILLER_44_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1144 U$$48/A1 U$$1174/A2 U$$50/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1145/A sky130_fd_sc_hd__a22o_1
XU$$1155 U$$1155/A U$$1163/B VGND VGND VPWR VPWR U$$1155/X sky130_fd_sc_hd__xor2_1
XU$$1166 U$$892/A1 U$$1194/A2 U$$894/A1 U$$1194/B2 VGND VGND VPWR VPWR U$$1167/A sky130_fd_sc_hd__a22o_1
XFILLER_31_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1177 U$$1177/A U$$1221/B VGND VGND VPWR VPWR U$$1177/X sky130_fd_sc_hd__xor2_1
XU$$1188 U$$503/A1 U$$1230/A2 U$$505/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1189/A sky130_fd_sc_hd__a22o_1
XU$$1199 U$$1199/A U$$1233/A VGND VGND VPWR VPWR U$$1199/X sky130_fd_sc_hd__xor2_1
XFILLER_148_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_111_0 dadda_fa_7_111_0/A dadda_fa_7_111_0/B dadda_fa_7_111_0/CIN VGND
+ VGND VPWR VPWR _408_/D _279_/D sky130_fd_sc_hd__fa_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_99_2 U$$3264/X U$$3397/X U$$3530/X VGND VGND VPWR VPWR dadda_fa_3_100_1/CIN
+ dadda_fa_3_99_3/B sky130_fd_sc_hd__fa_1
XFILLER_116_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_76_1 dadda_fa_5_76_1/A dadda_fa_5_76_1/B dadda_fa_5_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_77_0/B dadda_fa_7_76_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_69_0 dadda_fa_5_69_0/A dadda_fa_5_69_0/B dadda_fa_5_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_70_0/A dadda_fa_6_69_0/CIN sky130_fd_sc_hd__fa_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout707 U$$4190/B2 VGND VGND VPWR VPWR U$$4226/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout718 U$$3872/B2 VGND VGND VPWR VPWR U$$3892/B2 sky130_fd_sc_hd__buf_4
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout729 U$$3777/B2 VGND VGND VPWR VPWR U$$3773/B2 sky130_fd_sc_hd__buf_4
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_8 dadda_fa_1_68_8/A dadda_fa_1_68_8/B dadda_fa_1_68_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_69_3/A dadda_fa_3_68_0/A sky130_fd_sc_hd__fa_2
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_985 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3080 U$$3080/A1 U$$3124/A2 U$$4452/A1 U$$3124/B2 VGND VGND VPWR VPWR U$$3081/A
+ sky130_fd_sc_hd__a22o_1
XU$$3091 U$$3091/A U$$3151/A VGND VGND VPWR VPWR U$$3091/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_8_0 dadda_fa_6_8_0/A dadda_fa_6_8_0/B dadda_fa_6_8_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_9_0/B dadda_fa_7_8_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2390 U$$2390/A U$$2396/B VGND VGND VPWR VPWR U$$2390/X sky130_fd_sc_hd__xor2_1
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_71_0 dadda_fa_4_71_0/A dadda_fa_4_71_0/B dadda_fa_4_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_72_0/A dadda_fa_5_71_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_87_0 U$$1643/Y U$$1777/X U$$1910/X VGND VGND VPWR VPWR dadda_fa_2_88_3/A
+ dadda_fa_2_87_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$330 final_adder.U$$332/B final_adder.U$$330/B VGND VGND VPWR VPWR
+ final_adder.U$$456/B sky130_fd_sc_hd__and2_1
XFILLER_85_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$341 final_adder.U$$340/B final_adder.U$$215/X final_adder.U$$213/X
+ VGND VGND VPWR VPWR final_adder.U$$341/X sky130_fd_sc_hd__a21o_1
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$352 final_adder.U$$354/B final_adder.U$$352/B VGND VGND VPWR VPWR
+ final_adder.U$$478/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$363 final_adder.U$$362/B final_adder.U$$237/X final_adder.U$$235/X
+ VGND VGND VPWR VPWR final_adder.U$$363/X sky130_fd_sc_hd__a21o_1
XU$$202 U$$202/A U$$220/B VGND VGND VPWR VPWR U$$202/X sky130_fd_sc_hd__xor2_1
XFILLER_57_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$374 final_adder.U$$376/B final_adder.U$$374/B VGND VGND VPWR VPWR
+ final_adder.U$$500/B sky130_fd_sc_hd__and2_1
XFILLER_45_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$213 U$$76/A1 U$$213/A2 U$$78/A1 U$$213/B2 VGND VGND VPWR VPWR U$$214/A sky130_fd_sc_hd__a22o_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$385 final_adder.U$$384/B final_adder.U$$263/X final_adder.U$$259/X
+ VGND VGND VPWR VPWR final_adder.U$$385/X sky130_fd_sc_hd__a21o_1
XU$$224 U$$224/A U$$230/B VGND VGND VPWR VPWR U$$224/X sky130_fd_sc_hd__xor2_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$396 final_adder.U$$400/B final_adder.U$$396/B VGND VGND VPWR VPWR
+ final_adder.U$$520/B sky130_fd_sc_hd__and2_1
XU$$235 U$$370/B1 U$$271/A2 U$$922/A1 U$$271/B2 VGND VGND VPWR VPWR U$$236/A sky130_fd_sc_hd__a22o_1
XU$$246 U$$246/A U$$254/B VGND VGND VPWR VPWR U$$246/X sky130_fd_sc_hd__xor2_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$257 U$$805/A1 U$$271/A2 U$$805/B1 U$$271/B2 VGND VGND VPWR VPWR U$$258/A sky130_fd_sc_hd__a22o_1
XFILLER_72_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$268 U$$268/A U$$274/A VGND VGND VPWR VPWR U$$268/X sky130_fd_sc_hd__xor2_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$279 U$$277/B U$$273/A U$$275/A U$$274/Y VGND VGND VPWR VPWR U$$279/X sky130_fd_sc_hd__a22o_4
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$7 U$$7/A U$$9/B VGND VGND VPWR VPWR U$$7/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_86_0 dadda_fa_6_86_0/A dadda_fa_6_86_0/B dadda_fa_6_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_87_0/B dadda_fa_7_86_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_138_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$780 U$$780/A U$$820/B VGND VGND VPWR VPWR U$$780/X sky130_fd_sc_hd__xor2_1
XU$$791 U$$928/A1 U$$809/A2 U$$930/A1 U$$809/B2 VGND VGND VPWR VPWR U$$792/A sky130_fd_sc_hd__a22o_1
XFILLER_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_80_7 U$$3891/X U$$4024/X U$$4157/X VGND VGND VPWR VPWR dadda_fa_2_81_3/A
+ dadda_fa_2_80_5/CIN sky130_fd_sc_hd__fa_1
Xfanout504 U$$3245/A2 VGND VGND VPWR VPWR U$$3241/A2 sky130_fd_sc_hd__buf_4
XFILLER_59_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout515 U$$3018/X VGND VGND VPWR VPWR U$$3124/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_73_6 U$$4276/X U$$4409/X input227/X VGND VGND VPWR VPWR dadda_fa_2_74_2/B
+ dadda_fa_2_73_5/B sky130_fd_sc_hd__fa_1
Xfanout526 U$$3011/A2 VGND VGND VPWR VPWR U$$3005/A2 sky130_fd_sc_hd__buf_4
Xfanout537 U$$2844/A2 VGND VGND VPWR VPWR U$$2798/A2 sky130_fd_sc_hd__buf_4
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout548 U$$2607/X VGND VGND VPWR VPWR U$$2711/A2 sky130_fd_sc_hd__clkbuf_4
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout559 fanout561/X VGND VGND VPWR VPWR U$$2598/A2 sky130_fd_sc_hd__buf_6
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_66_5 input219/X dadda_fa_1_66_5/B dadda_fa_1_66_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_67_2/A dadda_fa_2_66_5/A sky130_fd_sc_hd__fa_1
XFILLER_112_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_59_4 U$$3184/X U$$3317/X U$$3450/X VGND VGND VPWR VPWR dadda_fa_2_60_1/CIN
+ dadda_fa_2_59_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1002 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_29_2 dadda_fa_4_29_2/A dadda_fa_4_29_2/B dadda_fa_4_29_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_30_0/CIN dadda_fa_5_29_1/CIN sky130_fd_sc_hd__fa_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4506 U$$4506/A1 U$$4388/X U$$4508/A1 U$$4506/B2 VGND VGND VPWR VPWR U$$4507/A
+ sky130_fd_sc_hd__a22o_1
XU$$4517 U$$4517/A U$$4517/B VGND VGND VPWR VPWR U$$4517/X sky130_fd_sc_hd__xor2_1
XFILLER_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3805 U$$4490/A1 U$$3833/A2 U$$4492/A1 U$$3833/B2 VGND VGND VPWR VPWR U$$3806/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_18_2 U$$841/X U$$974/X VGND VGND VPWR VPWR dadda_fa_4_19_1/CIN dadda_ha_3_18_2/SUM
+ sky130_fd_sc_hd__ha_1
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3816 U$$3816/A U$$3816/B VGND VGND VPWR VPWR U$$3816/X sky130_fd_sc_hd__xor2_1
XU$$3827 U$$4375/A1 U$$3829/A2 U$$4375/B1 U$$3829/B2 VGND VGND VPWR VPWR U$$3828/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$160 final_adder.U$$160/A final_adder.U$$160/B VGND VGND VPWR VPWR
+ final_adder.U$$288/B sky130_fd_sc_hd__and2_1
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3838 U$$3907/B VGND VGND VPWR VPWR U$$3838/Y sky130_fd_sc_hd__inv_1
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3849 U$$3849/A U$$3867/B VGND VGND VPWR VPWR U$$3849/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$171 final_adder.U$$170/B final_adder.U$$941/B1 final_adder.U$$171/B1
+ VGND VGND VPWR VPWR final_adder.U$$171/X sky130_fd_sc_hd__a21o_2
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$182 final_adder.U$$182/A final_adder.U$$182/B VGND VGND VPWR VPWR
+ final_adder.U$$310/B sky130_fd_sc_hd__and2_1
XFILLER_18_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_31_2 dadda_fa_3_31_2/A dadda_fa_3_31_2/B dadda_fa_3_31_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_32_1/A dadda_fa_4_31_2/B sky130_fd_sc_hd__fa_1
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$193 final_adder.U$$192/B final_adder.U$$963/B1 final_adder.U$$193/B1
+ VGND VGND VPWR VPWR final_adder.U$$193/X sky130_fd_sc_hd__a21o_1
XFILLER_46_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_24_1 U$$1119/X U$$1252/X U$$1385/X VGND VGND VPWR VPWR dadda_fa_4_25_0/CIN
+ dadda_fa_4_24_2/A sky130_fd_sc_hd__fa_1
XFILLER_73_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_17_0 U$$41/X U$$174/X U$$307/X VGND VGND VPWR VPWR dadda_fa_4_18_1/B dadda_fa_4_17_2/B
+ sky130_fd_sc_hd__fa_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_387_ _408_/CLK _387_/D VGND VGND VPWR VPWR _387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_83_5 dadda_fa_2_83_5/A dadda_fa_2_83_5/B dadda_fa_2_83_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_2/A dadda_fa_4_83_0/A sky130_fd_sc_hd__fa_2
XFILLER_114_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_76_4 dadda_fa_2_76_4/A dadda_fa_2_76_4/B dadda_fa_2_76_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_1/CIN dadda_fa_3_76_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_69_3 dadda_fa_2_69_3/A dadda_fa_2_69_3/B dadda_fa_2_69_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_1/B dadda_fa_3_69_3/B sky130_fd_sc_hd__fa_1
XFILLER_96_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_39_1 dadda_fa_5_39_1/A dadda_fa_5_39_1/B dadda_fa_5_39_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_40_0/B dadda_fa_7_39_0/A sky130_fd_sc_hd__fa_2
XFILLER_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_113_1 dadda_fa_5_113_1/A dadda_fa_5_113_1/B dadda_fa_5_113_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_114_0/B dadda_fa_7_113_0/A sky130_fd_sc_hd__fa_1
XFILLER_118_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_106_0 dadda_fa_5_106_0/A dadda_fa_5_106_0/B dadda_fa_5_106_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_107_0/A dadda_fa_6_106_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_71_3 U$$3341/X U$$3474/X U$$3607/X VGND VGND VPWR VPWR dadda_fa_2_72_1/B
+ dadda_fa_2_71_4/B sky130_fd_sc_hd__fa_1
XFILLER_114_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_2 U$$3327/X U$$3460/X U$$3593/X VGND VGND VPWR VPWR dadda_fa_2_65_1/A
+ dadda_fa_2_64_4/A sky130_fd_sc_hd__fa_1
XFILLER_59_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout389 U$$1087/A2 VGND VGND VPWR VPWR U$$981/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_4_41_1 dadda_fa_4_41_1/A dadda_fa_4_41_1/B dadda_fa_4_41_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_42_0/B dadda_fa_5_41_1/B sky130_fd_sc_hd__fa_1
XFILLER_100_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_57_1 U$$1584/X U$$1717/X U$$1850/X VGND VGND VPWR VPWR dadda_fa_2_58_0/CIN
+ dadda_fa_2_57_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_34_0 dadda_fa_4_34_0/A dadda_fa_4_34_0/B dadda_fa_4_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_35_0/A dadda_fa_5_34_1/A sky130_fd_sc_hd__fa_1
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ _328_/CLK _310_/D VGND VGND VPWR VPWR _310_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_241_ _377_/CLK _241_/D VGND VGND VPWR VPWR _241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_172_ _319_/CLK _172_/D VGND VGND VPWR VPWR _172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_86_3 dadda_fa_3_86_3/A dadda_fa_3_86_3/B dadda_fa_3_86_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_1/B dadda_fa_4_86_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_79_2 dadda_fa_3_79_2/A dadda_fa_3_79_2/B dadda_fa_3_79_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_1/A dadda_fa_4_79_2/B sky130_fd_sc_hd__fa_1
XFILLER_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_49_0 dadda_fa_6_49_0/A dadda_fa_6_49_0/B dadda_fa_6_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_50_0/B dadda_fa_7_49_0/CIN sky130_fd_sc_hd__fa_2
XU$$4303 U$$4440/A1 U$$4381/A2 U$$4440/B1 U$$4381/B2 VGND VGND VPWR VPWR U$$4304/A
+ sky130_fd_sc_hd__a22o_1
XU$$4314 U$$4314/A U$$4368/B VGND VGND VPWR VPWR U$$4314/X sky130_fd_sc_hd__xor2_1
XFILLER_120_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4325 U$$4460/B1 U$$4325/A2 U$$4464/A1 U$$4325/B2 VGND VGND VPWR VPWR U$$4326/A
+ sky130_fd_sc_hd__a22o_1
Xfanout890 U$$1480/B2 VGND VGND VPWR VPWR U$$1460/B2 sky130_fd_sc_hd__buf_4
XU$$4336 U$$4336/A U$$4350/B VGND VGND VPWR VPWR U$$4336/X sky130_fd_sc_hd__xor2_1
XU$$3602 U$$4287/A1 U$$3644/A2 U$$4426/A1 U$$3644/B2 VGND VGND VPWR VPWR U$$3603/A
+ sky130_fd_sc_hd__a22o_1
XU$$4347 U$$4482/B1 U$$4349/A2 U$$4349/A1 U$$4349/B2 VGND VGND VPWR VPWR U$$4348/A
+ sky130_fd_sc_hd__a22o_1
XU$$4358 U$$4358/A U$$4360/B VGND VGND VPWR VPWR U$$4358/X sky130_fd_sc_hd__xor2_1
XU$$3613 U$$3613/A U$$3659/B VGND VGND VPWR VPWR U$$3613/X sky130_fd_sc_hd__xor2_1
XU$$3624 U$$4309/A1 U$$3640/A2 U$$3763/A1 U$$3640/B2 VGND VGND VPWR VPWR U$$3625/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4369 U$$4506/A1 U$$4369/A2 U$$4508/A1 U$$4369/B2 VGND VGND VPWR VPWR U$$4370/A
+ sky130_fd_sc_hd__a22o_1
XU$$3635 U$$3635/A U$$3641/B VGND VGND VPWR VPWR U$$3635/X sky130_fd_sc_hd__xor2_1
XFILLER_133_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3646 U$$4468/A1 U$$3696/A2 U$$4470/A1 U$$3696/B2 VGND VGND VPWR VPWR U$$3647/A
+ sky130_fd_sc_hd__a22o_1
XU$$2901 U$$3447/B1 U$$2991/A2 U$$3314/A1 U$$2991/B2 VGND VGND VPWR VPWR U$$2902/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3657 U$$3657/A U$$3659/B VGND VGND VPWR VPWR U$$3657/X sky130_fd_sc_hd__xor2_1
XU$$2912 U$$2912/A U$$2990/B VGND VGND VPWR VPWR U$$2912/X sky130_fd_sc_hd__xor2_1
XU$$3668 U$$4214/B1 U$$3682/A2 U$$4492/A1 U$$3682/B2 VGND VGND VPWR VPWR U$$3669/A
+ sky130_fd_sc_hd__a22o_1
XU$$2923 U$$2923/A1 U$$2929/A2 U$$2925/A1 U$$2929/B2 VGND VGND VPWR VPWR U$$2924/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_108_2 dadda_fa_4_108_2/A dadda_fa_4_108_2/B dadda_fa_4_108_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_109_0/CIN dadda_fa_5_108_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2934 U$$2934/A U$$2938/B VGND VGND VPWR VPWR U$$2934/X sky130_fd_sc_hd__xor2_1
XU$$3679 U$$3679/A U$$3681/B VGND VGND VPWR VPWR U$$3679/X sky130_fd_sc_hd__xor2_1
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2945 U$$479/A1 U$$2989/A2 U$$479/B1 U$$2989/B2 VGND VGND VPWR VPWR U$$2946/A sky130_fd_sc_hd__a22o_1
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2956 U$$2956/A U$$2986/B VGND VGND VPWR VPWR U$$2956/X sky130_fd_sc_hd__xor2_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2967 U$$3239/B1 U$$2979/A2 U$$3106/A1 U$$2979/B2 VGND VGND VPWR VPWR U$$2968/A
+ sky130_fd_sc_hd__a22o_1
XU$$2978 U$$2978/A U$$3014/A VGND VGND VPWR VPWR U$$2978/X sky130_fd_sc_hd__xor2_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2989 U$$384/B1 U$$2989/A2 U$$251/A1 U$$2989/B2 VGND VGND VPWR VPWR U$$2990/A sky130_fd_sc_hd__a22o_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_892 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_81_2 dadda_fa_2_81_2/A dadda_fa_2_81_2/B dadda_fa_2_81_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_1/A dadda_fa_3_81_3/A sky130_fd_sc_hd__fa_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_74_1 dadda_fa_2_74_1/A dadda_fa_2_74_1/B dadda_fa_2_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_0/CIN dadda_fa_3_74_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_51_0 dadda_fa_5_51_0/A dadda_fa_5_51_0/B dadda_fa_5_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_52_0/A dadda_fa_6_51_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_2_67_0 dadda_fa_2_67_0/A dadda_fa_2_67_0/B dadda_fa_2_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_0/B dadda_fa_3_67_2/B sky130_fd_sc_hd__fa_1
XFILLER_96_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$907 final_adder.U$$136/A final_adder.U$$845/X final_adder.U$$907/B1
+ VGND VGND VPWR VPWR final_adder.U$$907/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$929 final_adder.U$$158/A final_adder.U$$867/X final_adder.U$$929/B1
+ VGND VGND VPWR VPWR final_adder.U$$929/X sky130_fd_sc_hd__a21o_1
XFILLER_68_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1044 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_clk _388_/CLK VGND VGND VPWR VPWR _384_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_96_2 dadda_fa_4_96_2/A dadda_fa_4_96_2/B dadda_fa_4_96_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_97_0/CIN dadda_fa_5_96_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_89_1 dadda_fa_4_89_1/A dadda_fa_4_89_1/B dadda_fa_4_89_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_90_0/B dadda_fa_5_89_1/B sky130_fd_sc_hd__fa_1
XFILLER_106_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_66_0 dadda_fa_7_66_0/A dadda_fa_7_66_0/B dadda_fa_7_66_0/CIN VGND VGND
+ VPWR VPWR _363_/D _234_/D sky130_fd_sc_hd__fa_1
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1107 U$$3751/B1 VGND VGND VPWR VPWR U$$4162/B1 sky130_fd_sc_hd__buf_6
XFILLER_154_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1118 U$$3338/A1 VGND VGND VPWR VPWR U$$596/B1 sky130_fd_sc_hd__buf_4
Xfanout1129 U$$870/A1 VGND VGND VPWR VPWR U$$48/A1 sky130_fd_sc_hd__buf_4
XFILLER_102_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2208 U$$973/B1 U$$2252/A2 U$$840/A1 U$$2252/B2 VGND VGND VPWR VPWR U$$2209/A sky130_fd_sc_hd__a22o_1
XU$$2219 U$$2219/A U$$2231/B VGND VGND VPWR VPWR U$$2219/X sky130_fd_sc_hd__xor2_1
XFILLER_27_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1507 U$$1507/A VGND VGND VPWR VPWR U$$1507/Y sky130_fd_sc_hd__inv_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1518 U$$1518/A U$$1568/B VGND VGND VPWR VPWR U$$1518/X sky130_fd_sc_hd__xor2_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1529 U$$2625/A1 U$$1567/A2 U$$983/A1 U$$1567/B2 VGND VGND VPWR VPWR U$$1530/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_clk _370_/CLK VGND VGND VPWR VPWR _377_/CLK sky130_fd_sc_hd__clkbuf_16
X_224_ _356_/CLK _224_/D VGND VGND VPWR VPWR _224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_91_1 dadda_fa_3_91_1/A dadda_fa_3_91_1/B dadda_fa_3_91_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_0/CIN dadda_fa_4_91_2/A sky130_fd_sc_hd__fa_1
XFILLER_171_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_84_0 dadda_fa_3_84_0/A dadda_fa_3_84_0/B dadda_fa_3_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_0/B dadda_fa_4_84_1/CIN sky130_fd_sc_hd__fa_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4253_1835 VGND VGND VPWR VPWR U$$4253_1835/HI U$$4253/A1 sky130_fd_sc_hd__conb_1
XFILLER_111_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1630 input115/X VGND VGND VPWR VPWR U$$940/A1 sky130_fd_sc_hd__buf_4
XFILLER_66_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1641 input114/X VGND VGND VPWR VPWR U$$251/B1 sky130_fd_sc_hd__buf_2
XU$$4100 U$$4100/A U$$4108/B VGND VGND VPWR VPWR U$$4100/X sky130_fd_sc_hd__xor2_1
Xfanout1652 U$$4498/A1 VGND VGND VPWR VPWR U$$4359/B1 sky130_fd_sc_hd__buf_2
XFILLER_78_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4111 input57/X VGND VGND VPWR VPWR U$$4113/B sky130_fd_sc_hd__inv_1
Xfanout1663 input112/X VGND VGND VPWR VPWR U$$2578/A1 sky130_fd_sc_hd__buf_8
XU$$4122 U$$4257/B1 U$$4158/A2 U$$4259/B1 U$$4158/B2 VGND VGND VPWR VPWR U$$4123/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1674 U$$2711/A1 VGND VGND VPWR VPWR U$$930/A1 sky130_fd_sc_hd__buf_4
XU$$4133 U$$4133/A U$$4133/B VGND VGND VPWR VPWR U$$4133/X sky130_fd_sc_hd__xor2_1
Xfanout1685 U$$1320/B VGND VGND VPWR VPWR U$$1282/B sky130_fd_sc_hd__buf_6
XFILLER_93_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4144 U$$4416/B1 U$$4190/A2 U$$4283/A1 U$$4190/B2 VGND VGND VPWR VPWR U$$4145/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1696 U$$975/A1 VGND VGND VPWR VPWR U$$16/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_168_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4155 U$$4155/A U$$4175/B VGND VGND VPWR VPWR U$$4155/X sky130_fd_sc_hd__xor2_1
XU$$3410 U$$3684/A1 U$$3418/A2 U$$3684/B1 U$$3418/B2 VGND VGND VPWR VPWR U$$3411/A
+ sky130_fd_sc_hd__a22o_1
XU$$4166 U$$4440/A1 U$$4174/A2 U$$4440/B1 U$$4174/B2 VGND VGND VPWR VPWR U$$4167/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_46_5 dadda_fa_2_46_5/A dadda_fa_2_46_5/B dadda_fa_2_46_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_2/A dadda_fa_4_46_0/A sky130_fd_sc_hd__fa_1
XU$$3421 U$$3421/A U$$3424/A VGND VGND VPWR VPWR U$$3421/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_113_0 U$$4223/X U$$4356/X U$$4489/X VGND VGND VPWR VPWR dadda_fa_5_114_0/A
+ dadda_fa_5_113_1/A sky130_fd_sc_hd__fa_1
XFILLER_19_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4177 U$$4177/A U$$4247/A VGND VGND VPWR VPWR U$$4177/X sky130_fd_sc_hd__xor2_1
XU$$3432 U$$3432/A U$$3468/B VGND VGND VPWR VPWR U$$3432/X sky130_fd_sc_hd__xor2_1
XFILLER_65_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4188 U$$4460/B1 U$$4190/A2 U$$4464/A1 U$$4190/B2 VGND VGND VPWR VPWR U$$4189/A
+ sky130_fd_sc_hd__a22o_1
XU$$3443 U$$3580/A1 U$$3523/A2 U$$3580/B1 U$$3523/B2 VGND VGND VPWR VPWR U$$3444/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3454 U$$3454/A U$$3468/B VGND VGND VPWR VPWR U$$3454/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_39_4 input189/X dadda_fa_2_39_4/B dadda_fa_2_39_4/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_40_1/CIN dadda_fa_3_39_3/CIN sky130_fd_sc_hd__fa_1
XU$$4199 U$$4199/A U$$4215/B VGND VGND VPWR VPWR U$$4199/X sky130_fd_sc_hd__xor2_1
XU$$3465 U$$4287/A1 U$$3505/A2 U$$4426/A1 U$$3505/B2 VGND VGND VPWR VPWR U$$3466/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2720 U$$2720/A U$$2739/A VGND VGND VPWR VPWR U$$2720/X sky130_fd_sc_hd__xor2_1
XU$$2731 U$$3416/A1 U$$2737/A2 U$$3418/A1 U$$2737/B2 VGND VGND VPWR VPWR U$$2732/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3476 U$$3476/A U$$3482/B VGND VGND VPWR VPWR U$$3476/X sky130_fd_sc_hd__xor2_1
XU$$2742 U$$2841/B VGND VGND VPWR VPWR U$$2742/Y sky130_fd_sc_hd__inv_1
XU$$3487 U$$4307/B1 U$$3511/A2 U$$3763/A1 U$$3511/B2 VGND VGND VPWR VPWR U$$3488/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2753 U$$2753/A U$$2799/B VGND VGND VPWR VPWR U$$2753/X sky130_fd_sc_hd__xor2_1
XU$$3498 U$$3498/A U$$3506/B VGND VGND VPWR VPWR U$$3498/X sky130_fd_sc_hd__xor2_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2764 U$$981/B1 U$$2804/A2 U$$985/A1 U$$2804/B2 VGND VGND VPWR VPWR U$$2765/A sky130_fd_sc_hd__a22o_1
XU$$2775 U$$2775/A U$$2811/B VGND VGND VPWR VPWR U$$2775/X sky130_fd_sc_hd__xor2_1
XU$$2786 U$$2923/A1 U$$2804/A2 U$$2925/A1 U$$2804/B2 VGND VGND VPWR VPWR U$$2787/A
+ sky130_fd_sc_hd__a22o_1
XU$$2797 U$$2797/A U$$2841/B VGND VGND VPWR VPWR U$$2797/X sky130_fd_sc_hd__xor2_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_13_clk _370_/CLK VGND VGND VPWR VPWR _397_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_99_0 dadda_fa_5_99_0/A dadda_fa_5_99_0/B dadda_fa_5_99_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_100_0/A dadda_fa_6_99_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$704 final_adder.U$$720/B final_adder.U$$704/B VGND VGND VPWR VPWR
+ final_adder.U$$784/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$715 final_adder.U$$714/B final_adder.U$$611/X final_adder.U$$595/X
+ VGND VGND VPWR VPWR final_adder.U$$715/X sky130_fd_sc_hd__a21o_1
XFILLER_68_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$737 final_adder.U$$720/A final_adder.U$$255/X final_adder.U$$617/X
+ VGND VGND VPWR VPWR final_adder.U$$737/X sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$748 final_adder.U$$780/B final_adder.U$$748/B VGND VGND VPWR VPWR
+ final_adder.U$$748/X sky130_fd_sc_hd__and2_1
XFILLER_112_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$759 final_adder.U$$758/B final_adder.U$$679/X final_adder.U$$647/X
+ VGND VGND VPWR VPWR final_adder.U$$759/X sky130_fd_sc_hd__a21o_1
XU$$609 U$$609/A U$$643/B VGND VGND VPWR VPWR U$$609/X sky130_fd_sc_hd__xor2_1
XFILLER_71_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_108_1 U$$3681/X U$$3814/X U$$3947/X VGND VGND VPWR VPWR dadda_fa_4_109_0/CIN
+ dadda_fa_4_108_2/A sky130_fd_sc_hd__fa_1
XFILLER_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput290 output290/A VGND VGND VPWR VPWR o[14] sky130_fd_sc_hd__buf_2
XFILLER_0_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_49_3 dadda_fa_3_49_3/A dadda_fa_3_49_3/B dadda_fa_3_49_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_1/B dadda_fa_4_49_2/CIN sky130_fd_sc_hd__fa_1
XU$$2005 U$$2005/A U$$2031/B VGND VGND VPWR VPWR U$$2005/X sky130_fd_sc_hd__xor2_1
XFILLER_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2016 U$$920/A1 U$$2052/A2 U$$920/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2017/A sky130_fd_sc_hd__a22o_1
XU$$2027 U$$2027/A U$$2043/B VGND VGND VPWR VPWR U$$2027/X sky130_fd_sc_hd__xor2_1
XU$$2038 U$$2312/A1 U$$2044/A2 U$$2175/B1 U$$2044/B2 VGND VGND VPWR VPWR U$$2039/A
+ sky130_fd_sc_hd__a22o_1
XU$$1304 U$$1304/A U$$1320/B VGND VGND VPWR VPWR U$$1304/X sky130_fd_sc_hd__xor2_1
XU$$2049 U$$2049/A U$$2053/B VGND VGND VPWR VPWR U$$2049/X sky130_fd_sc_hd__xor2_1
XFILLER_43_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1315 U$$82/A1 U$$1353/A2 U$$3920/A1 U$$1353/B2 VGND VGND VPWR VPWR U$$1316/A sky130_fd_sc_hd__a22o_1
XU$$1326 U$$1326/A U$$1328/B VGND VGND VPWR VPWR U$$1326/X sky130_fd_sc_hd__xor2_1
XU$$1337 U$$926/A1 U$$1361/A2 U$$928/A1 U$$1361/B2 VGND VGND VPWR VPWR U$$1338/A sky130_fd_sc_hd__a22o_1
XU$$1348 U$$1348/A U$$1358/B VGND VGND VPWR VPWR U$$1348/X sky130_fd_sc_hd__xor2_1
XFILLER_128_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1359 U$$811/A1 U$$1359/A2 U$$811/B1 U$$1359/B2 VGND VGND VPWR VPWR U$$1360/A sky130_fd_sc_hd__a22o_1
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_207_ _344_/CLK _207_/D VGND VGND VPWR VPWR _207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_954 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1120 final_adder.U$$158/A final_adder.U$$867/X VGND VGND VPWR VPWR
+ output380/A sky130_fd_sc_hd__xor2_1
XFILLER_128_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1131 final_adder.U$$148/B final_adder.U$$919/X VGND VGND VPWR VPWR
+ output265/A sky130_fd_sc_hd__xor2_1
XFILLER_172_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1142 final_adder.U$$136/A final_adder.U$$845/X VGND VGND VPWR VPWR
+ output277/A sky130_fd_sc_hd__xor2_1
XFILLER_156_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_clk _201_/CLK VGND VGND VPWR VPWR _319_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_931 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1460 U$$2015/B VGND VGND VPWR VPWR U$$1971/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_51_3 dadda_fa_2_51_3/A dadda_fa_2_51_3/B dadda_fa_2_51_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_1/B dadda_fa_3_51_3/B sky130_fd_sc_hd__fa_1
XU$$4411_1853 VGND VGND VPWR VPWR U$$4411_1853/HI U$$4411/B sky130_fd_sc_hd__conb_1
XFILLER_39_858 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1471 U$$1882/B VGND VGND VPWR VPWR U$$1854/B sky130_fd_sc_hd__buf_6
Xfanout1482 U$$1741/B VGND VGND VPWR VPWR U$$1777/B sky130_fd_sc_hd__clkbuf_8
Xfanout1493 U$$1608/B VGND VGND VPWR VPWR U$$1630/B sky130_fd_sc_hd__clkbuf_4
XFILLER_65_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_44_2 U$$3061/B input195/X dadda_fa_2_44_2/CIN VGND VGND VPWR VPWR dadda_fa_3_45_1/A
+ dadda_fa_3_44_3/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$11 _307_/Q _179_/Q VGND VGND VPWR VPWR final_adder.U$$245/B1 final_adder.U$$244/B
+ sky130_fd_sc_hd__ha_1
XFILLER_38_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3240 U$$3240/A U$$3242/B VGND VGND VPWR VPWR U$$3240/X sky130_fd_sc_hd__xor2_1
XFILLER_80_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_21_1 dadda_fa_5_21_1/A dadda_fa_5_21_1/B dadda_fa_5_21_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_22_0/B dadda_fa_7_21_0/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$22 _318_/Q _190_/Q VGND VGND VPWR VPWR final_adder.U$$233/A2 final_adder.U$$232/A
+ sky130_fd_sc_hd__ha_1
XU$$3251 U$$4482/B1 U$$3251/A2 U$$4349/A1 U$$3251/B2 VGND VGND VPWR VPWR U$$3252/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$33 _329_/Q _201_/Q VGND VGND VPWR VPWR final_adder.U$$223/B1 final_adder.U$$222/B
+ sky130_fd_sc_hd__ha_1
XU$$3262 U$$3262/A U$$3284/B VGND VGND VPWR VPWR U$$3262/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_37_1 U$$1145/X U$$1278/X U$$1411/X VGND VGND VPWR VPWR dadda_fa_3_38_0/CIN
+ dadda_fa_3_37_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$44 _340_/Q _212_/Q VGND VGND VPWR VPWR final_adder.U$$981/B1 final_adder.U$$210/A
+ sky130_fd_sc_hd__ha_1
XFILLER_94_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3273 U$$4093/B1 U$$3285/A2 U$$3960/A1 U$$3285/B2 VGND VGND VPWR VPWR U$$3274/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$55 _351_/Q _223_/Q VGND VGND VPWR VPWR final_adder.U$$201/B1 final_adder.U$$200/B
+ sky130_fd_sc_hd__ha_1
XFILLER_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$66 _362_/Q _234_/Q VGND VGND VPWR VPWR final_adder.U$$959/B1 final_adder.U$$188/A
+ sky130_fd_sc_hd__ha_2
XU$$3284 U$$3284/A U$$3284/B VGND VGND VPWR VPWR U$$3284/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_14_0 dadda_fa_5_14_0/A dadda_fa_5_14_0/B dadda_fa_5_14_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_15_0/A dadda_fa_6_14_0/CIN sky130_fd_sc_hd__fa_1
XU$$3295 U$$3295/A U$$3335/B VGND VGND VPWR VPWR U$$3295/X sky130_fd_sc_hd__xor2_1
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2550 U$$4331/A1 U$$2600/A2 U$$4196/A1 U$$2600/B2 VGND VGND VPWR VPWR U$$2551/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$77 _373_/Q _245_/Q VGND VGND VPWR VPWR final_adder.U$$179/B1 final_adder.U$$178/B
+ sky130_fd_sc_hd__ha_1
XU$$2561 U$$2561/A U$$2603/A VGND VGND VPWR VPWR U$$2561/X sky130_fd_sc_hd__xor2_1
XFILLER_80_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2572 U$$2707/B1 U$$2574/A2 U$$2574/A1 U$$2574/B2 VGND VGND VPWR VPWR U$$2573/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$88 _384_/Q _256_/Q VGND VGND VPWR VPWR final_adder.U$$937/B1 final_adder.U$$166/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$99 _395_/Q _267_/Q VGND VGND VPWR VPWR final_adder.U$$157/B1 final_adder.U$$156/B
+ sky130_fd_sc_hd__ha_1
XFILLER_80_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2583 U$$2583/A U$$2591/B VGND VGND VPWR VPWR U$$2583/X sky130_fd_sc_hd__xor2_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2594 U$$950/A1 U$$2600/A2 U$$952/A1 U$$2600/B2 VGND VGND VPWR VPWR U$$2595/A sky130_fd_sc_hd__a22o_1
XFILLER_61_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1860 U$$1860/A U$$1882/B VGND VGND VPWR VPWR U$$1860/X sky130_fd_sc_hd__xor2_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1871 U$$88/B1 U$$1909/A2 U$$503/A1 U$$1909/B2 VGND VGND VPWR VPWR U$$1872/A sky130_fd_sc_hd__a22o_1
XU$$1882 U$$1882/A U$$1882/B VGND VGND VPWR VPWR U$$1882/X sky130_fd_sc_hd__xor2_1
XFILLER_166_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1893 U$$2576/B1 U$$1911/A2 U$$388/A1 U$$1911/B2 VGND VGND VPWR VPWR U$$1894/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_40_3 U$$1284/X U$$1417/X VGND VGND VPWR VPWR dadda_fa_2_41_4/CIN dadda_fa_3_40_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_130_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_59_2 dadda_fa_4_59_2/A dadda_fa_4_59_2/B dadda_fa_4_59_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_60_0/CIN dadda_fa_5_59_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$501 final_adder.U$$500/B final_adder.U$$379/X final_adder.U$$375/X
+ VGND VGND VPWR VPWR final_adder.U$$501/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$512 final_adder.U$$520/B final_adder.U$$512/B VGND VGND VPWR VPWR
+ final_adder.U$$632/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$523 final_adder.U$$522/B final_adder.U$$407/X final_adder.U$$399/X
+ VGND VGND VPWR VPWR final_adder.U$$523/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$534 final_adder.U$$542/B final_adder.U$$534/B VGND VGND VPWR VPWR
+ final_adder.U$$654/B sky130_fd_sc_hd__and2_1
Xdadda_ha_4_10_1 U$$426/X U$$559/X VGND VGND VPWR VPWR dadda_fa_5_11_1/A dadda_ha_4_10_1/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_56_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$545 final_adder.U$$544/B final_adder.U$$429/X final_adder.U$$421/X
+ VGND VGND VPWR VPWR final_adder.U$$545/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$556 final_adder.U$$564/B final_adder.U$$556/B VGND VGND VPWR VPWR
+ final_adder.U$$676/B sky130_fd_sc_hd__and2_1
Xdadda_fa_7_29_0 dadda_fa_7_29_0/A dadda_fa_7_29_0/B dadda_fa_7_29_0/CIN VGND VGND
+ VPWR VPWR _326_/D _197_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$567 final_adder.U$$566/B final_adder.U$$451/X final_adder.U$$443/X
+ VGND VGND VPWR VPWR final_adder.U$$567/X sky130_fd_sc_hd__a21o_1
XU$$406 U$$406/A1 U$$406/A2 U$$406/B1 U$$406/B2 VGND VGND VPWR VPWR U$$407/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$578 final_adder.U$$586/B final_adder.U$$578/B VGND VGND VPWR VPWR
+ final_adder.U$$698/B sky130_fd_sc_hd__and2_1
XFILLER_45_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$417 U$$417/A1 U$$447/A2 U$$965/B1 U$$447/B2 VGND VGND VPWR VPWR U$$418/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$589 final_adder.U$$588/B final_adder.U$$473/X final_adder.U$$465/X
+ VGND VGND VPWR VPWR final_adder.U$$589/X sky130_fd_sc_hd__a21o_1
XU$$428 U$$428/A U$$480/B VGND VGND VPWR VPWR U$$428/X sky130_fd_sc_hd__xor2_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$439 U$$576/A1 U$$505/A2 U$$576/B1 U$$505/B2 VGND VGND VPWR VPWR U$$440/A sky130_fd_sc_hd__a22o_1
XFILLER_72_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_61_2 dadda_fa_3_61_2/A dadda_fa_3_61_2/B dadda_fa_3_61_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_1/A dadda_fa_4_61_2/B sky130_fd_sc_hd__fa_1
XFILLER_94_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_54_1 dadda_fa_3_54_1/A dadda_fa_3_54_1/B dadda_fa_3_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_0/CIN dadda_fa_4_54_2/A sky130_fd_sc_hd__fa_1
XFILLER_85_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_31_0 dadda_fa_6_31_0/A dadda_fa_6_31_0/B dadda_fa_6_31_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_32_0/B dadda_fa_7_31_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_87_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_47_0 dadda_fa_3_47_0/A dadda_fa_3_47_0/B dadda_fa_3_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_0/B dadda_fa_4_47_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$940 U$$940/A1 U$$942/A2 U$$942/A1 U$$942/B2 VGND VGND VPWR VPWR U$$941/A sky130_fd_sc_hd__a22o_1
XFILLER_62_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$951 U$$951/A U$$958/A VGND VGND VPWR VPWR U$$951/X sky130_fd_sc_hd__xor2_1
XU$$1101 U$$1099/B U$$962/A input8/X U$$1096/Y VGND VGND VPWR VPWR U$$1101/X sky130_fd_sc_hd__a22o_1
XU$$962 U$$962/A U$$962/B VGND VGND VPWR VPWR U$$962/X sky130_fd_sc_hd__and2_1
XFILLER_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$973 U$$973/A1 U$$979/A2 U$$973/B1 U$$979/B2 VGND VGND VPWR VPWR U$$974/A sky130_fd_sc_hd__a22o_1
XU$$1112 U$$16/A1 U$$1174/A2 U$$18/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1113/A sky130_fd_sc_hd__a22o_1
XU$$1123 U$$1123/A U$$1163/B VGND VGND VPWR VPWR U$$1123/X sky130_fd_sc_hd__xor2_1
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$984 U$$984/A U$$998/B VGND VGND VPWR VPWR U$$984/X sky130_fd_sc_hd__xor2_1
XU$$995 U$$995/A1 U$$997/A2 U$$997/A1 U$$997/B2 VGND VGND VPWR VPWR U$$996/A sky130_fd_sc_hd__a22o_1
XU$$1134 U$$721/B1 U$$1170/A2 U$$999/A1 U$$1170/B2 VGND VGND VPWR VPWR U$$1135/A sky130_fd_sc_hd__a22o_1
XU$$1145 U$$1145/A U$$1175/B VGND VGND VPWR VPWR U$$1145/X sky130_fd_sc_hd__xor2_1
XFILLER_16_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1156 U$$60/A1 U$$1164/A2 U$$62/A1 U$$1164/B2 VGND VGND VPWR VPWR U$$1157/A sky130_fd_sc_hd__a22o_1
XU$$1167 U$$1167/A U$$1189/B VGND VGND VPWR VPWR U$$1167/X sky130_fd_sc_hd__xor2_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1178 U$$82/A1 U$$1218/A2 U$$82/B1 U$$1218/B2 VGND VGND VPWR VPWR U$$1179/A sky130_fd_sc_hd__a22o_1
XFILLER_31_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1189 U$$1189/A U$$1189/B VGND VGND VPWR VPWR U$$1189/X sky130_fd_sc_hd__xor2_1
XU$$4441_1868 VGND VGND VPWR VPWR U$$4441_1868/HI U$$4441/B sky130_fd_sc_hd__conb_1
XFILLER_8_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_104_0 dadda_fa_7_104_0/A dadda_fa_7_104_0/B dadda_fa_7_104_0/CIN VGND
+ VGND VPWR VPWR _401_/D _272_/D sky130_fd_sc_hd__fa_1
XFILLER_129_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4517_1906 VGND VGND VPWR VPWR U$$4517_1906/HI U$$4517/B sky130_fd_sc_hd__conb_1
XFILLER_102_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_99_3 U$$3663/X U$$3796/X U$$3929/X VGND VGND VPWR VPWR dadda_fa_3_100_2/A
+ dadda_fa_3_99_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_98_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_5_69_1 dadda_fa_5_69_1/A dadda_fa_5_69_1/B dadda_fa_5_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_70_0/B dadda_fa_7_69_0/A sky130_fd_sc_hd__fa_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout708 U$$4115/X VGND VGND VPWR VPWR U$$4190/B2 sky130_fd_sc_hd__buf_6
XFILLER_59_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout719 U$$3912/B2 VGND VGND VPWR VPWR U$$3872/B2 sky130_fd_sc_hd__clkbuf_4
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1290 fanout1299/X VGND VGND VPWR VPWR U$$4026/B sky130_fd_sc_hd__buf_6
XFILLER_67_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3070 U$$4027/B1 U$$3072/A2 U$$4442/A1 U$$3072/B2 VGND VGND VPWR VPWR U$$3071/A
+ sky130_fd_sc_hd__a22o_1
XU$$3081 U$$3081/A U$$3123/B VGND VGND VPWR VPWR U$$3081/X sky130_fd_sc_hd__xor2_1
XU$$3092 U$$3638/B1 U$$3108/A2 U$$3503/B1 U$$3108/B2 VGND VGND VPWR VPWR U$$3093/A
+ sky130_fd_sc_hd__a22o_1
XU$$2380 U$$2380/A U$$2416/B VGND VGND VPWR VPWR U$$2380/X sky130_fd_sc_hd__xor2_1
XU$$2391 U$$2665/A1 U$$2395/A2 U$$2665/B1 U$$2395/B2 VGND VGND VPWR VPWR U$$2392/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1690 U$$729/B1 U$$1696/A2 U$$596/A1 U$$1696/B2 VGND VGND VPWR VPWR U$$1691/A sky130_fd_sc_hd__a22o_1
XFILLER_136_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_71_1 dadda_fa_4_71_1/A dadda_fa_4_71_1/B dadda_fa_4_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_72_0/B dadda_fa_5_71_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_87_1 U$$2043/X U$$2176/X U$$2309/X VGND VGND VPWR VPWR dadda_fa_2_88_3/B
+ dadda_fa_2_87_5/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_64_0 dadda_fa_4_64_0/A dadda_fa_4_64_0/B dadda_fa_4_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_65_0/A dadda_fa_5_64_1/A sky130_fd_sc_hd__fa_1
XFILLER_131_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$320 final_adder.U$$322/B final_adder.U$$320/B VGND VGND VPWR VPWR
+ final_adder.U$$446/B sky130_fd_sc_hd__and2_1
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$331 final_adder.U$$330/B final_adder.U$$205/X final_adder.U$$203/X
+ VGND VGND VPWR VPWR final_adder.U$$331/X sky130_fd_sc_hd__a21o_1
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$342 final_adder.U$$344/B final_adder.U$$342/B VGND VGND VPWR VPWR
+ final_adder.U$$468/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$353 final_adder.U$$352/B final_adder.U$$227/X final_adder.U$$225/X
+ VGND VGND VPWR VPWR final_adder.U$$353/X sky130_fd_sc_hd__a21o_1
XFILLER_85_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$364 final_adder.U$$366/B final_adder.U$$364/B VGND VGND VPWR VPWR
+ final_adder.U$$490/B sky130_fd_sc_hd__and2_1
XU$$203 U$$66/A1 U$$219/A2 U$$66/B1 U$$219/B2 VGND VGND VPWR VPWR U$$204/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$375 final_adder.U$$374/B final_adder.U$$249/X final_adder.U$$247/X
+ VGND VGND VPWR VPWR final_adder.U$$375/X sky130_fd_sc_hd__a21o_1
XFILLER_57_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$214 U$$214/A U$$214/B VGND VGND VPWR VPWR U$$214/X sky130_fd_sc_hd__xor2_1
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$386 final_adder.U$$390/B final_adder.U$$386/B VGND VGND VPWR VPWR
+ final_adder.U$$510/B sky130_fd_sc_hd__and2_1
XU$$225 U$$499/A1 U$$229/A2 U$$90/A1 U$$229/B2 VGND VGND VPWR VPWR U$$226/A sky130_fd_sc_hd__a22o_1
XFILLER_45_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$397 final_adder.U$$396/B final_adder.U$$275/X final_adder.U$$271/X
+ VGND VGND VPWR VPWR final_adder.U$$397/X sky130_fd_sc_hd__a21o_1
XU$$236 U$$236/A U$$273/A VGND VGND VPWR VPWR U$$236/X sky130_fd_sc_hd__xor2_1
XFILLER_72_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$247 U$$384/A1 U$$253/A2 U$$384/B1 U$$253/B2 VGND VGND VPWR VPWR U$$248/A sky130_fd_sc_hd__a22o_1
XFILLER_33_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$258 U$$258/A U$$274/A VGND VGND VPWR VPWR U$$258/X sky130_fd_sc_hd__xor2_1
XU$$269 U$$406/A1 U$$271/A2 U$$406/B1 U$$271/B2 VGND VGND VPWR VPWR U$$270/A sky130_fd_sc_hd__a22o_1
XFILLER_72_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$8 U$$8/A1 U$$8/A2 U$$8/B1 U$$8/B2 VGND VGND VPWR VPWR U$$9/A sky130_fd_sc_hd__a22o_1
XFILLER_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_76_1 U$$1223/X U$$1356/X VGND VGND VPWR VPWR dadda_fa_1_77_8/CIN dadda_fa_2_76_0/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_6_79_0 dadda_fa_6_79_0/A dadda_fa_6_79_0/B dadda_fa_6_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_80_0/B dadda_fa_7_79_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$770 U$$770/A U$$821/A VGND VGND VPWR VPWR U$$770/X sky130_fd_sc_hd__xor2_1
XU$$781 U$$781/A1 U$$817/A2 U$$783/A1 U$$817/B2 VGND VGND VPWR VPWR U$$782/A sky130_fd_sc_hd__a22o_1
XU$$792 U$$792/A U$$804/B VGND VGND VPWR VPWR U$$792/X sky130_fd_sc_hd__xor2_1
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_81_0 dadda_fa_5_81_0/A dadda_fa_5_81_0/B dadda_fa_5_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_82_0/A dadda_fa_6_81_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_97_0 U$$2328/Y U$$2462/X U$$2595/X VGND VGND VPWR VPWR dadda_fa_3_98_0/B
+ dadda_fa_3_97_2/B sky130_fd_sc_hd__fa_1
XFILLER_6_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout505 U$$3155/X VGND VGND VPWR VPWR U$$3245/A2 sky130_fd_sc_hd__buf_2
Xfanout516 U$$3018/X VGND VGND VPWR VPWR U$$3122/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout527 U$$2881/X VGND VGND VPWR VPWR U$$3011/A2 sky130_fd_sc_hd__buf_4
Xfanout538 U$$2844/A2 VGND VGND VPWR VPWR U$$2804/A2 sky130_fd_sc_hd__buf_4
XFILLER_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_73_7 dadda_fa_1_73_7/A dadda_fa_1_73_7/B dadda_fa_1_73_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_74_2/CIN dadda_fa_2_73_5/CIN sky130_fd_sc_hd__fa_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout549 U$$2679/A2 VGND VGND VPWR VPWR U$$2681/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_82_0_1924 VGND VGND VPWR VPWR dadda_fa_1_82_0/A dadda_fa_1_82_0_1924/LO
+ sky130_fd_sc_hd__conb_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_66_6 dadda_fa_1_66_6/A dadda_fa_1_66_6/B dadda_fa_1_66_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_67_2/B dadda_fa_2_66_5/B sky130_fd_sc_hd__fa_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_59_5 U$$3583/X U$$3716/X U$$3849/X VGND VGND VPWR VPWR dadda_fa_2_60_2/A
+ dadda_fa_2_59_5/A sky130_fd_sc_hd__fa_1
XFILLER_132_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_96_0 dadda_fa_7_96_0/A dadda_fa_7_96_0/B dadda_fa_7_96_0/CIN VGND VGND
+ VPWR VPWR _393_/D _264_/D sky130_fd_sc_hd__fa_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4507 U$$4507/A U$$4507/B VGND VGND VPWR VPWR U$$4507/X sky130_fd_sc_hd__xor2_1
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_111_0 dadda_fa_6_111_0/A dadda_fa_6_111_0/B dadda_fa_6_111_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_112_0/B dadda_fa_7_111_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3806 U$$3806/A U$$3835/A VGND VGND VPWR VPWR U$$3806/X sky130_fd_sc_hd__xor2_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3817 U$$3817/A1 U$$3829/A2 U$$3817/B1 U$$3829/B2 VGND VGND VPWR VPWR U$$3818/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$150 final_adder.U$$150/A final_adder.U$$150/B VGND VGND VPWR VPWR
+ final_adder.U$$278/B sky130_fd_sc_hd__and2_1
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3828 U$$3828/A U$$3828/B VGND VGND VPWR VPWR U$$3828/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$161 final_adder.U$$160/B final_adder.U$$931/B1 final_adder.U$$161/B1
+ VGND VGND VPWR VPWR final_adder.U$$161/X sky130_fd_sc_hd__a21o_1
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$172 final_adder.U$$172/A final_adder.U$$172/B VGND VGND VPWR VPWR
+ final_adder.U$$300/B sky130_fd_sc_hd__and2_1
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3839 U$$3973/A U$$3839/B VGND VGND VPWR VPWR U$$3839/X sky130_fd_sc_hd__and2_1
Xdadda_fa_3_31_3 dadda_fa_3_31_3/A dadda_fa_3_31_3/B dadda_fa_3_31_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_32_1/B dadda_fa_4_31_2/CIN sky130_fd_sc_hd__fa_1
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$183 final_adder.U$$182/B final_adder.U$$953/B1 final_adder.U$$183/B1
+ VGND VGND VPWR VPWR final_adder.U$$183/X sky130_fd_sc_hd__a21o_1
XFILLER_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$194 final_adder.U$$194/A final_adder.U$$194/B VGND VGND VPWR VPWR
+ final_adder.U$$322/B sky130_fd_sc_hd__and2_1
XFILLER_18_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_24_2 U$$1518/X U$$1651/X U$$1699/B VGND VGND VPWR VPWR dadda_fa_4_25_1/A
+ dadda_fa_4_24_2/B sky130_fd_sc_hd__fa_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_386_ _386_/CLK _386_/D VGND VGND VPWR VPWR _386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_76_5 dadda_fa_2_76_5/A dadda_fa_2_76_5/B dadda_fa_2_76_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_2/A dadda_fa_4_76_0/A sky130_fd_sc_hd__fa_2
XFILLER_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_69_4 dadda_fa_2_69_4/A dadda_fa_2_69_4/B dadda_fa_2_69_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_1/CIN dadda_fa_3_69_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_150_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput190 c[3] VGND VGND VPWR VPWR input190/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_106_1 dadda_fa_5_106_1/A dadda_fa_5_106_1/B dadda_fa_5_106_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_107_0/B dadda_fa_7_106_0/A sky130_fd_sc_hd__fa_1
XFILLER_117_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4493_1894 VGND VGND VPWR VPWR U$$4493_1894/HI U$$4493/B sky130_fd_sc_hd__conb_1
XFILLER_160_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_71_4 U$$3740/X U$$3873/X U$$4006/X VGND VGND VPWR VPWR dadda_fa_2_72_1/CIN
+ dadda_fa_2_71_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_64_3 U$$3726/X U$$3859/X U$$3992/X VGND VGND VPWR VPWR dadda_fa_2_65_1/B
+ dadda_fa_2_64_4/B sky130_fd_sc_hd__fa_1
XFILLER_100_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_41_2 dadda_fa_4_41_2/A dadda_fa_4_41_2/B dadda_fa_4_41_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_42_0/CIN dadda_fa_5_41_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_57_2 U$$1983/X U$$2116/X U$$2249/X VGND VGND VPWR VPWR dadda_fa_2_58_1/A
+ dadda_fa_2_57_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_34_1 dadda_fa_4_34_1/A dadda_fa_4_34_1/B dadda_fa_4_34_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_35_0/B dadda_fa_5_34_1/B sky130_fd_sc_hd__fa_1
XFILLER_27_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_11_0 dadda_fa_7_11_0/A dadda_fa_7_11_0/B dadda_fa_7_11_0/CIN VGND VGND
+ VPWR VPWR _308_/D _179_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_27_0 dadda_fa_4_27_0/A dadda_fa_4_27_0/B dadda_fa_4_27_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_28_0/A dadda_fa_5_27_1/A sky130_fd_sc_hd__fa_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_240_ _369_/CLK _240_/D VGND VGND VPWR VPWR _240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_171_ _319_/CLK _171_/D VGND VGND VPWR VPWR _171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_0_60_4 U$$1723/X U$$1856/X VGND VGND VPWR VPWR dadda_fa_1_61_7/B dadda_fa_2_60_0/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_3_79_3 dadda_fa_3_79_3/A dadda_fa_3_79_3/B dadda_fa_3_79_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_1/B dadda_fa_4_79_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4304 U$$4304/A U$$4384/A VGND VGND VPWR VPWR U$$4304/X sky130_fd_sc_hd__xor2_1
XU$$4315 U$$4315/A1 U$$4373/A2 U$$4315/B1 U$$4373/B2 VGND VGND VPWR VPWR U$$4316/A
+ sky130_fd_sc_hd__a22o_1
Xfanout880 U$$259/B2 VGND VGND VPWR VPWR U$$229/B2 sky130_fd_sc_hd__buf_4
XU$$4326 U$$4326/A U$$4350/B VGND VGND VPWR VPWR U$$4326/X sky130_fd_sc_hd__xor2_1
XFILLER_77_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout891 U$$1452/B2 VGND VGND VPWR VPWR U$$1414/B2 sky130_fd_sc_hd__buf_4
XU$$4337 U$$4474/A1 U$$4359/A2 U$$4474/B1 U$$4359/B2 VGND VGND VPWR VPWR U$$4338/A
+ sky130_fd_sc_hd__a22o_1
XU$$3603 U$$3603/A U$$3607/B VGND VGND VPWR VPWR U$$3603/X sky130_fd_sc_hd__xor2_1
XU$$4348 U$$4348/A U$$4350/B VGND VGND VPWR VPWR U$$4348/X sky130_fd_sc_hd__xor2_1
XFILLER_46_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3614 U$$3751/A1 U$$3656/A2 U$$3751/B1 U$$3656/B2 VGND VGND VPWR VPWR U$$3615/A
+ sky130_fd_sc_hd__a22o_1
XU$$4359 U$$4359/A1 U$$4359/A2 U$$4359/B1 U$$4359/B2 VGND VGND VPWR VPWR U$$4360/A
+ sky130_fd_sc_hd__a22o_1
XU$$3625 U$$3625/A U$$3641/B VGND VGND VPWR VPWR U$$3625/X sky130_fd_sc_hd__xor2_1
XU$$3636 U$$3908/B1 U$$3640/A2 U$$3636/B1 U$$3640/B2 VGND VGND VPWR VPWR U$$3637/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3647 U$$3647/A U$$3695/B VGND VGND VPWR VPWR U$$3647/X sky130_fd_sc_hd__xor2_1
XU$$2902 U$$2902/A U$$2944/B VGND VGND VPWR VPWR U$$2902/X sky130_fd_sc_hd__xor2_1
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2913 U$$3048/B1 U$$2991/A2 U$$4011/A1 U$$2991/B2 VGND VGND VPWR VPWR U$$2914/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3658 U$$4478/B1 U$$3658/A2 U$$4345/A1 U$$3658/B2 VGND VGND VPWR VPWR U$$3659/A
+ sky130_fd_sc_hd__a22o_1
XU$$3669 U$$3669/A U$$3681/B VGND VGND VPWR VPWR U$$3669/X sky130_fd_sc_hd__xor2_1
XU$$2924 U$$2924/A U$$2926/B VGND VGND VPWR VPWR U$$2924/X sky130_fd_sc_hd__xor2_1
XFILLER_46_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2935 U$$4442/A1 U$$2937/A2 U$$4442/B1 U$$2937/B2 VGND VGND VPWR VPWR U$$2936/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2946 U$$2946/A U$$2990/B VGND VGND VPWR VPWR U$$2946/X sky130_fd_sc_hd__xor2_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2957 U$$3642/A1 U$$2979/A2 U$$3642/B1 U$$2979/B2 VGND VGND VPWR VPWR U$$2958/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2968 U$$2968/A U$$2974/B VGND VGND VPWR VPWR U$$2968/X sky130_fd_sc_hd__xor2_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2979 U$$922/B1 U$$2979/A2 U$$2979/B1 U$$2979/B2 VGND VGND VPWR VPWR U$$2980/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_369_ _369_/CLK _369_/D VGND VGND VPWR VPWR _369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_81_3 dadda_fa_2_81_3/A dadda_fa_2_81_3/B dadda_fa_2_81_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_1/B dadda_fa_3_81_3/B sky130_fd_sc_hd__fa_1
XFILLER_114_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_74_2 dadda_fa_2_74_2/A dadda_fa_2_74_2/B dadda_fa_2_74_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_1/A dadda_fa_3_74_3/A sky130_fd_sc_hd__fa_1
XFILLER_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_51_1 dadda_fa_5_51_1/A dadda_fa_5_51_1/B dadda_fa_5_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_52_0/B dadda_fa_7_51_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_67_1 dadda_fa_2_67_1/A dadda_fa_2_67_1/B dadda_fa_2_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_0/CIN dadda_fa_3_67_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_867 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_44_0 dadda_fa_5_44_0/A dadda_fa_5_44_0/B dadda_fa_5_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_45_0/A dadda_fa_6_44_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$919 final_adder.U$$148/A final_adder.U$$857/X final_adder.U$$919/B1
+ VGND VGND VPWR VPWR final_adder.U$$919/X sky130_fd_sc_hd__a21o_1
XFILLER_3_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_89_2 dadda_fa_4_89_2/A dadda_fa_4_89_2/B dadda_fa_4_89_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_90_0/CIN dadda_fa_5_89_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_133_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_59_0 dadda_fa_7_59_0/A dadda_fa_7_59_0/B dadda_fa_7_59_0/CIN VGND VGND
+ VPWR VPWR _356_/D _227_/D sky130_fd_sc_hd__fa_1
XFILLER_161_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1108 U$$3751/B1 VGND VGND VPWR VPWR U$$4438/A1 sky130_fd_sc_hd__buf_2
XFILLER_99_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1119 U$$3338/A1 VGND VGND VPWR VPWR U$$735/A1 sky130_fd_sc_hd__buf_4
XFILLER_87_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_62_0 U$$2392/X U$$2525/X U$$2658/X VGND VGND VPWR VPWR dadda_fa_2_63_0/B
+ dadda_fa_2_62_3/B sky130_fd_sc_hd__fa_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2209 U$$2209/A U$$2253/B VGND VGND VPWR VPWR U$$2209/X sky130_fd_sc_hd__xor2_1
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1508 input15/X VGND VGND VPWR VPWR U$$1510/B sky130_fd_sc_hd__inv_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1519 U$$2887/B1 U$$1567/A2 U$$2754/A1 U$$1567/B2 VGND VGND VPWR VPWR U$$1520/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_223_ _353_/CLK _223_/D VGND VGND VPWR VPWR _223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_91_2 dadda_fa_3_91_2/A dadda_fa_3_91_2/B dadda_fa_3_91_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_1/A dadda_fa_4_91_2/B sky130_fd_sc_hd__fa_1
XFILLER_109_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_84_1 dadda_fa_3_84_1/A dadda_fa_3_84_1/B dadda_fa_3_84_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_0/CIN dadda_fa_4_84_2/A sky130_fd_sc_hd__fa_1
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_61_0 dadda_fa_6_61_0/A dadda_fa_6_61_0/B dadda_fa_6_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_62_0/B dadda_fa_7_61_0/CIN sky130_fd_sc_hd__fa_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_77_0 dadda_fa_3_77_0/A dadda_fa_3_77_0/B dadda_fa_3_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_0/B dadda_fa_4_77_1/CIN sky130_fd_sc_hd__fa_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1620 input116/X VGND VGND VPWR VPWR U$$942/A1 sky130_fd_sc_hd__buf_6
XFILLER_111_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1631 U$$2993/B1 VGND VGND VPWR VPWR U$$253/B1 sky130_fd_sc_hd__buf_6
Xfanout1642 U$$4500/A1 VGND VGND VPWR VPWR U$$4363/A1 sky130_fd_sc_hd__buf_4
Xfanout1653 U$$2578/B1 VGND VGND VPWR VPWR U$$4498/A1 sky130_fd_sc_hd__clkbuf_4
XU$$4101 U$$4375/A1 U$$4105/A2 U$$4375/B1 U$$4105/B2 VGND VGND VPWR VPWR U$$4102/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1664 U$$2711/B1 VGND VGND VPWR VPWR U$$932/A1 sky130_fd_sc_hd__buf_4
XU$$4112 U$$4247/A VGND VGND VPWR VPWR U$$4112/Y sky130_fd_sc_hd__inv_1
XU$$4123 U$$4123/A U$$4133/B VGND VGND VPWR VPWR U$$4123/X sky130_fd_sc_hd__xor2_1
Xfanout1675 fanout1680/X VGND VGND VPWR VPWR U$$654/B1 sky130_fd_sc_hd__clkbuf_8
XU$$4134 U$$4271/A1 U$$4244/A2 U$$985/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4135/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1686 U$$1320/B VGND VGND VPWR VPWR U$$1278/B sky130_fd_sc_hd__clkbuf_4
XU$$3400 U$$3948/A1 U$$3416/A2 U$$3948/B1 U$$3416/B2 VGND VGND VPWR VPWR U$$3401/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1697 U$$562/B1 VGND VGND VPWR VPWR U$$975/A1 sky130_fd_sc_hd__buf_2
XU$$4145 U$$4145/A U$$4191/B VGND VGND VPWR VPWR U$$4145/X sky130_fd_sc_hd__xor2_1
XU$$4156 U$$4430/A1 U$$4174/A2 U$$4158/A1 U$$4174/B2 VGND VGND VPWR VPWR U$$4157/A
+ sky130_fd_sc_hd__a22o_1
XU$$3411 U$$3411/A U$$3411/B VGND VGND VPWR VPWR U$$3411/X sky130_fd_sc_hd__xor2_1
XU$$3422 U$$4107/A1 U$$3422/A2 U$$3422/B1 U$$3422/B2 VGND VGND VPWR VPWR U$$3423/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_113_1 input144/X dadda_fa_4_113_1/B dadda_fa_4_113_1/CIN VGND VGND VPWR
+ VPWR dadda_fa_5_114_0/B dadda_fa_5_113_1/B sky130_fd_sc_hd__fa_1
XU$$4167 U$$4167/A U$$4175/B VGND VGND VPWR VPWR U$$4167/X sky130_fd_sc_hd__xor2_1
XFILLER_19_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3433 U$$3981/A1 U$$3473/A2 U$$4257/A1 U$$3473/B2 VGND VGND VPWR VPWR U$$3434/A
+ sky130_fd_sc_hd__a22o_1
XU$$4178 U$$4315/A1 U$$4240/A2 U$$4454/A1 U$$4240/B2 VGND VGND VPWR VPWR U$$4179/A
+ sky130_fd_sc_hd__a22o_1
XU$$4189 U$$4189/A U$$4191/B VGND VGND VPWR VPWR U$$4189/X sky130_fd_sc_hd__xor2_1
XU$$3444 U$$3444/A U$$3482/B VGND VGND VPWR VPWR U$$3444/X sky130_fd_sc_hd__xor2_1
XFILLER_34_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3455 U$$4001/B1 U$$3471/A2 U$$854/A1 U$$3471/B2 VGND VGND VPWR VPWR U$$3456/A
+ sky130_fd_sc_hd__a22o_1
XU$$2710 U$$2710/A U$$2740/A VGND VGND VPWR VPWR U$$2710/X sky130_fd_sc_hd__xor2_1
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3466 U$$3466/A U$$3506/B VGND VGND VPWR VPWR U$$3466/X sky130_fd_sc_hd__xor2_1
XFILLER_74_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_39_5 dadda_fa_2_39_5/A dadda_fa_2_39_5/B dadda_fa_2_39_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_40_2/A dadda_fa_4_39_0/A sky130_fd_sc_hd__fa_1
XFILLER_92_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2721 U$$3817/A1 U$$2737/A2 U$$120/A1 U$$2737/B2 VGND VGND VPWR VPWR U$$2722/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_106_0 dadda_fa_4_106_0/A dadda_fa_4_106_0/B dadda_fa_4_106_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_107_0/A dadda_fa_5_106_1/A sky130_fd_sc_hd__fa_1
XU$$2732 U$$2732/A U$$2738/B VGND VGND VPWR VPWR U$$2732/X sky130_fd_sc_hd__xor2_1
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3477 input79/X U$$3523/A2 U$$876/A1 U$$3523/B2 VGND VGND VPWR VPWR U$$3478/A sky130_fd_sc_hd__a22o_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2743 U$$2877/A U$$2743/B VGND VGND VPWR VPWR U$$2743/X sky130_fd_sc_hd__and2_1
XU$$3488 U$$3488/A U$$3562/A VGND VGND VPWR VPWR U$$3488/X sky130_fd_sc_hd__xor2_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2754 U$$2754/A1 U$$2798/A2 U$$2891/B1 U$$2798/B2 VGND VGND VPWR VPWR U$$2755/A
+ sky130_fd_sc_hd__a22o_1
XU$$3499 U$$3499/A1 U$$3505/A2 U$$3636/B1 U$$3505/B2 VGND VGND VPWR VPWR U$$3500/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2765 U$$2765/A U$$2805/B VGND VGND VPWR VPWR U$$2765/X sky130_fd_sc_hd__xor2_1
XU$$2776 U$$4283/A1 U$$2856/A2 U$$4011/A1 U$$2856/B2 VGND VGND VPWR VPWR U$$2777/A
+ sky130_fd_sc_hd__a22o_1
XU$$2787 U$$2787/A U$$2805/B VGND VGND VPWR VPWR U$$2787/X sky130_fd_sc_hd__xor2_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2798 U$$4442/A1 U$$2798/A2 U$$4442/B1 U$$2798/B2 VGND VGND VPWR VPWR U$$2799/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_99_1 dadda_fa_5_99_1/A dadda_fa_5_99_1/B dadda_fa_5_99_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_100_0/B dadda_fa_7_99_0/A sky130_fd_sc_hd__fa_1
XFILLER_147_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$705 final_adder.U$$704/B final_adder.U$$601/X final_adder.U$$585/X
+ VGND VGND VPWR VPWR final_adder.U$$705/X sky130_fd_sc_hd__a21o_1
XFILLER_84_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$716 final_adder.U$$716/A final_adder.U$$716/B VGND VGND VPWR VPWR
+ final_adder.U$$796/A sky130_fd_sc_hd__and2_1
XFILLER_57_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$727 final_adder.U$$710/A final_adder.U$$623/X final_adder.U$$607/X
+ VGND VGND VPWR VPWR final_adder.U$$727/X sky130_fd_sc_hd__a21o_2
XFILLER_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$749 final_adder.U$$748/B final_adder.U$$669/X final_adder.U$$637/X
+ VGND VGND VPWR VPWR final_adder.U$$749/X sky130_fd_sc_hd__a21o_1
XFILLER_110_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_94_0 dadda_fa_4_94_0/A dadda_fa_4_94_0/B dadda_fa_4_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_95_0/A dadda_fa_5_94_1/A sky130_fd_sc_hd__fa_1
XFILLER_4_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_108_2 U$$4080/X U$$4213/X U$$4346/X VGND VGND VPWR VPWR dadda_fa_4_109_1/A
+ dadda_fa_4_108_2/B sky130_fd_sc_hd__fa_1
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput280 output280/A VGND VGND VPWR VPWR o[120] sky130_fd_sc_hd__buf_2
XFILLER_88_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput291 output291/A VGND VGND VPWR VPWR o[15] sky130_fd_sc_hd__buf_2
XFILLER_59_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2006 U$$88/A1 U$$2006/A2 U$$88/B1 U$$2006/B2 VGND VGND VPWR VPWR U$$2007/A sky130_fd_sc_hd__a22o_1
XFILLER_56_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2017 U$$2017/A U$$2053/B VGND VGND VPWR VPWR U$$2017/X sky130_fd_sc_hd__xor2_1
XU$$2028 U$$2576/A1 U$$2044/A2 U$$2576/B1 U$$2044/B2 VGND VGND VPWR VPWR U$$2029/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2039 U$$2039/A U$$2043/B VGND VGND VPWR VPWR U$$2039/X sky130_fd_sc_hd__xor2_1
XFILLER_74_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1305 U$$72/A1 U$$1309/A2 U$$74/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1306/A sky130_fd_sc_hd__a22o_1
XU$$1316 U$$1316/A U$$1320/B VGND VGND VPWR VPWR U$$1316/X sky130_fd_sc_hd__xor2_1
XU$$1327 U$$94/A1 U$$1327/A2 U$$96/A1 U$$1327/B2 VGND VGND VPWR VPWR U$$1328/A sky130_fd_sc_hd__a22o_1
XFILLER_71_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1338 U$$1338/A U$$1364/B VGND VGND VPWR VPWR U$$1338/X sky130_fd_sc_hd__xor2_1
XU$$1349 U$$253/A1 U$$1359/A2 U$$253/B1 U$$1359/B2 VGND VGND VPWR VPWR U$$1350/A sky130_fd_sc_hd__a22o_1
XFILLER_129_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_206_ _353_/CLK _206_/D VGND VGND VPWR VPWR _206_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$1110 final_adder.U$$168/A final_adder.U$$877/X VGND VGND VPWR VPWR
+ output369/A sky130_fd_sc_hd__xor2_1
XFILLER_128_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1121 final_adder.U$$158/B final_adder.U$$929/X VGND VGND VPWR VPWR
+ output381/A sky130_fd_sc_hd__xor2_1
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1132 final_adder.U$$146/A final_adder.U$$855/X VGND VGND VPWR VPWR
+ output266/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1143 final_adder.U$$136/B final_adder.U$$907/X VGND VGND VPWR VPWR
+ output278/A sky130_fd_sc_hd__xor2_1
XFILLER_156_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1450 U$$2140/B VGND VGND VPWR VPWR U$$2130/B sky130_fd_sc_hd__buf_8
Xfanout1461 U$$2015/B VGND VGND VPWR VPWR U$$1981/B sky130_fd_sc_hd__clkbuf_4
Xfanout1472 input20/X VGND VGND VPWR VPWR U$$1882/B sky130_fd_sc_hd__buf_6
XFILLER_94_943 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_51_4 dadda_fa_2_51_4/A dadda_fa_2_51_4/B dadda_fa_2_51_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_1/CIN dadda_fa_3_51_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1483 U$$1781/A VGND VGND VPWR VPWR U$$1741/B sky130_fd_sc_hd__buf_6
Xfanout1494 U$$1626/B VGND VGND VPWR VPWR U$$1608/B sky130_fd_sc_hd__buf_6
XFILLER_65_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_44_3 dadda_fa_2_44_3/A dadda_fa_2_44_3/B dadda_fa_2_44_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_45_1/B dadda_fa_3_44_3/B sky130_fd_sc_hd__fa_1
XU$$3230 U$$3230/A U$$3242/B VGND VGND VPWR VPWR U$$3230/X sky130_fd_sc_hd__xor2_1
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$12 _308_/Q _180_/Q VGND VGND VPWR VPWR final_adder.U$$243/A2 final_adder.U$$242/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3241 U$$3376/B1 U$$3241/A2 U$$3243/A1 U$$3241/B2 VGND VGND VPWR VPWR U$$3242/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$23 _319_/Q _191_/Q VGND VGND VPWR VPWR final_adder.U$$233/B1 final_adder.U$$232/B
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$34 _330_/Q _202_/Q VGND VGND VPWR VPWR final_adder.U$$991/B1 final_adder.U$$220/A
+ sky130_fd_sc_hd__ha_1
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_37_2 U$$1544/X U$$1677/X U$$1810/X VGND VGND VPWR VPWR dadda_fa_3_38_1/A
+ dadda_fa_3_37_3/A sky130_fd_sc_hd__fa_1
XU$$3252 U$$3252/A U$$3287/A VGND VGND VPWR VPWR U$$3252/X sky130_fd_sc_hd__xor2_1
XU$$3263 U$$3948/A1 U$$3283/A2 U$$3948/B1 U$$3283/B2 VGND VGND VPWR VPWR U$$3264/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$45 _341_/Q _213_/Q VGND VGND VPWR VPWR final_adder.U$$211/B1 final_adder.U$$210/B
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3274 U$$3274/A U$$3286/B VGND VGND VPWR VPWR U$$3274/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$56 _352_/Q _224_/Q VGND VGND VPWR VPWR final_adder.U$$969/B1 final_adder.U$$198/A
+ sky130_fd_sc_hd__ha_1
XU$$2540 U$$2814/A1 U$$2540/A2 U$$74/B1 U$$2540/B2 VGND VGND VPWR VPWR U$$2541/A sky130_fd_sc_hd__a22o_1
XFILLER_94_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3285 U$$3285/A1 U$$3285/A2 U$$3285/B1 U$$3285/B2 VGND VGND VPWR VPWR U$$3286/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$67 _363_/Q _235_/Q VGND VGND VPWR VPWR final_adder.U$$189/B1 final_adder.U$$188/B
+ sky130_fd_sc_hd__ha_2
XU$$2551 U$$2551/A U$$2591/B VGND VGND VPWR VPWR U$$2551/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_14_1 dadda_fa_5_14_1/A dadda_fa_5_14_1/B dadda_fa_5_14_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_15_0/B dadda_fa_7_14_0/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$78 _374_/Q _246_/Q VGND VGND VPWR VPWR final_adder.U$$947/B1 final_adder.U$$176/A
+ sky130_fd_sc_hd__ha_1
XU$$3296 U$$4392/A1 U$$3338/A2 U$$3296/B1 U$$3338/B2 VGND VGND VPWR VPWR U$$3297/A
+ sky130_fd_sc_hd__a22o_1
XU$$2562 U$$2973/A1 U$$2574/A2 U$$2973/B1 U$$2574/B2 VGND VGND VPWR VPWR U$$2563/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2573 U$$2573/A U$$2575/B VGND VGND VPWR VPWR U$$2573/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$89 _385_/Q _257_/Q VGND VGND VPWR VPWR final_adder.U$$167/B1 final_adder.U$$166/B
+ sky130_fd_sc_hd__ha_4
XU$$2584 U$$4365/A1 U$$2598/A2 U$$4365/B1 U$$2598/B2 VGND VGND VPWR VPWR U$$2585/A
+ sky130_fd_sc_hd__a22o_1
XU$$2595 U$$2595/A U$$2602/A VGND VGND VPWR VPWR U$$2595/X sky130_fd_sc_hd__xor2_1
XU$$1850 U$$1850/A U$$1854/B VGND VGND VPWR VPWR U$$1850/X sky130_fd_sc_hd__xor2_1
XU$$1861 U$$3503/B1 U$$1909/A2 U$$3370/A1 U$$1909/B2 VGND VGND VPWR VPWR U$$1862/A
+ sky130_fd_sc_hd__a22o_1
XU$$1872 U$$1872/A U$$1874/B VGND VGND VPWR VPWR U$$1872/X sky130_fd_sc_hd__xor2_1
XFILLER_61_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1883 U$$787/A1 U$$1915/A2 U$$787/B1 U$$1915/B2 VGND VGND VPWR VPWR U$$1884/A sky130_fd_sc_hd__a22o_1
XU$$1894 U$$1894/A U$$1910/B VGND VGND VPWR VPWR U$$1894/X sky130_fd_sc_hd__xor2_1
XFILLER_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_945 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$513 final_adder.U$$512/B final_adder.U$$397/X final_adder.U$$389/X
+ VGND VGND VPWR VPWR final_adder.U$$513/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$524 final_adder.U$$532/B final_adder.U$$524/B VGND VGND VPWR VPWR
+ final_adder.U$$644/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$535 final_adder.U$$534/B final_adder.U$$419/X final_adder.U$$411/X
+ VGND VGND VPWR VPWR final_adder.U$$535/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$546 final_adder.U$$554/B final_adder.U$$546/B VGND VGND VPWR VPWR
+ final_adder.U$$666/B sky130_fd_sc_hd__and2_1
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$557 final_adder.U$$556/B final_adder.U$$441/X final_adder.U$$433/X
+ VGND VGND VPWR VPWR final_adder.U$$557/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$568 final_adder.U$$576/B final_adder.U$$568/B VGND VGND VPWR VPWR
+ final_adder.U$$688/B sky130_fd_sc_hd__and2_1
XU$$407 U$$407/A U$$407/B VGND VGND VPWR VPWR U$$407/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$579 final_adder.U$$578/B final_adder.U$$463/X final_adder.U$$455/X
+ VGND VGND VPWR VPWR final_adder.U$$579/X sky130_fd_sc_hd__a21o_1
XU$$418 U$$418/A U$$448/B VGND VGND VPWR VPWR U$$418/X sky130_fd_sc_hd__xor2_1
XFILLER_38_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$429 U$$566/A1 U$$447/A2 U$$979/A1 U$$447/B2 VGND VGND VPWR VPWR U$$430/A sky130_fd_sc_hd__a22o_1
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4427_1861 VGND VGND VPWR VPWR U$$4427_1861/HI U$$4427/B sky130_fd_sc_hd__conb_1
XFILLER_53_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_113_0 U$$3424/Y U$$3558/X U$$3691/X VGND VGND VPWR VPWR dadda_fa_4_114_1/CIN
+ dadda_fa_4_113_2/B sky130_fd_sc_hd__fa_1
XFILLER_109_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_61_3 dadda_fa_3_61_3/A dadda_fa_3_61_3/B dadda_fa_3_61_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_1/B dadda_fa_4_61_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$828_1914 VGND VGND VPWR VPWR U$$828_1914/HI U$$828/A1 sky130_fd_sc_hd__conb_1
Xdadda_fa_3_54_2 dadda_fa_3_54_2/A dadda_fa_3_54_2/B dadda_fa_3_54_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_1/A dadda_fa_4_54_2/B sky130_fd_sc_hd__fa_1
XFILLER_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_47_1 dadda_fa_3_47_1/A dadda_fa_3_47_1/B dadda_fa_3_47_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_0/CIN dadda_fa_4_47_2/A sky130_fd_sc_hd__fa_1
XFILLER_91_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_24_0 dadda_fa_6_24_0/A dadda_fa_6_24_0/B dadda_fa_6_24_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_25_0/B dadda_fa_7_24_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_90_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$930 U$$930/A1 U$$942/A2 U$$932/A1 U$$942/B2 VGND VGND VPWR VPWR U$$931/A sky130_fd_sc_hd__a22o_1
XU$$941 U$$941/A U$$943/B VGND VGND VPWR VPWR U$$941/X sky130_fd_sc_hd__xor2_1
XFILLER_165_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$952 U$$952/A1 U$$952/A2 U$$954/A1 U$$952/B2 VGND VGND VPWR VPWR U$$953/A sky130_fd_sc_hd__a22o_1
XU$$963 U$$961/Y input6/X U$$959/A U$$962/X U$$959/Y VGND VGND VPWR VPWR U$$963/X
+ sky130_fd_sc_hd__a32o_4
XU$$1102 U$$1102/A1 U$$1170/A2 U$$967/A1 U$$1170/B2 VGND VGND VPWR VPWR U$$1103/A
+ sky130_fd_sc_hd__a22o_1
XU$$974 U$$974/A U$$980/B VGND VGND VPWR VPWR U$$974/X sky130_fd_sc_hd__xor2_1
XU$$1113 U$$1113/A U$$1175/B VGND VGND VPWR VPWR U$$1113/X sky130_fd_sc_hd__xor2_1
XU$$1124 U$$850/A1 U$$1164/A2 U$$989/A1 U$$1164/B2 VGND VGND VPWR VPWR U$$1125/A sky130_fd_sc_hd__a22o_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$985 U$$985/A1 U$$999/A2 U$$987/A1 U$$999/B2 VGND VGND VPWR VPWR U$$986/A sky130_fd_sc_hd__a22o_1
XU$$996 U$$996/A U$$998/B VGND VGND VPWR VPWR U$$996/X sky130_fd_sc_hd__xor2_1
XU$$1135 U$$1135/A U$$1171/B VGND VGND VPWR VPWR U$$1135/X sky130_fd_sc_hd__xor2_1
XU$$1146 U$$50/A1 U$$1170/A2 U$$50/B1 U$$1170/B2 VGND VGND VPWR VPWR U$$1147/A sky130_fd_sc_hd__a22o_1
XU$$1157 U$$1157/A U$$1163/B VGND VGND VPWR VPWR U$$1157/X sky130_fd_sc_hd__xor2_1
XFILLER_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1168 U$$894/A1 U$$1202/A2 U$$896/A1 U$$1202/B2 VGND VGND VPWR VPWR U$$1169/A sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_112_2 U$$4088/X U$$4221/X VGND VGND VPWR VPWR dadda_fa_4_113_2/A dadda_ha_3_112_2/SUM
+ sky130_fd_sc_hd__ha_1
XU$$1179 U$$1179/A U$$1221/B VGND VGND VPWR VPWR U$$1179/X sky130_fd_sc_hd__xor2_1
XFILLER_129_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_99_4 U$$4062/X U$$4195/X U$$4328/X VGND VGND VPWR VPWR dadda_fa_3_100_2/B
+ dadda_fa_4_99_0/A sky130_fd_sc_hd__fa_2
XFILLER_132_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout709 U$$4043/B2 VGND VGND VPWR VPWR U$$4025/B2 sky130_fd_sc_hd__clkbuf_4
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1280 input56/X VGND VGND VPWR VPWR U$$363/B sky130_fd_sc_hd__buf_6
XFILLER_67_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1291 fanout1299/X VGND VGND VPWR VPWR U$$4006/B sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_2_42_0 U$$1953/X U$$2086/X U$$2219/X VGND VGND VPWR VPWR dadda_fa_3_43_0/B
+ dadda_fa_3_42_2/B sky130_fd_sc_hd__fa_1
XFILLER_93_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3060 U$$4430/A1 U$$3072/A2 U$$4158/A1 U$$3072/B2 VGND VGND VPWR VPWR U$$3061/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3071 U$$3071/A U$$3073/B VGND VGND VPWR VPWR U$$3071/X sky130_fd_sc_hd__xor2_1
XU$$3082 U$$4315/A1 U$$3118/A2 U$$4454/A1 U$$3118/B2 VGND VGND VPWR VPWR U$$3083/A
+ sky130_fd_sc_hd__a22o_1
XU$$3093 U$$3093/A U$$3107/B VGND VGND VPWR VPWR U$$3093/X sky130_fd_sc_hd__xor2_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2370 U$$2370/A U$$2412/B VGND VGND VPWR VPWR U$$2370/X sky130_fd_sc_hd__xor2_1
XFILLER_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2381 U$$874/A1 U$$2415/A2 U$$876/A1 U$$2415/B2 VGND VGND VPWR VPWR U$$2382/A sky130_fd_sc_hd__a22o_1
XU$$2392 U$$2392/A U$$2396/B VGND VGND VPWR VPWR U$$2392/X sky130_fd_sc_hd__xor2_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1680 U$$36/A1 U$$1702/A2 U$$38/A1 U$$1702/B2 VGND VGND VPWR VPWR U$$1681/A sky130_fd_sc_hd__a22o_1
XU$$1691 U$$1691/A U$$1697/B VGND VGND VPWR VPWR U$$1691/X sky130_fd_sc_hd__xor2_1
XFILLER_139_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_88_4 U$$3242/X U$$3375/X VGND VGND VPWR VPWR dadda_fa_2_89_4/CIN dadda_fa_3_88_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_136_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4457_1876 VGND VGND VPWR VPWR U$$4457_1876/HI U$$4457/B sky130_fd_sc_hd__conb_1
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_71_2 dadda_fa_4_71_2/A dadda_fa_4_71_2/B dadda_fa_4_71_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_72_0/CIN dadda_fa_5_71_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_162_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_87_2 U$$2442/X U$$2575/X U$$2708/X VGND VGND VPWR VPWR dadda_fa_2_88_3/CIN
+ dadda_fa_2_87_5/B sky130_fd_sc_hd__fa_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_64_1 dadda_fa_4_64_1/A dadda_fa_4_64_1/B dadda_fa_4_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_65_0/B dadda_fa_5_64_1/B sky130_fd_sc_hd__fa_1
XFILLER_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_41_0 dadda_fa_7_41_0/A dadda_fa_7_41_0/B dadda_fa_7_41_0/CIN VGND VGND
+ VPWR VPWR _338_/D _209_/D sky130_fd_sc_hd__fa_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_57_0 dadda_fa_4_57_0/A dadda_fa_4_57_0/B dadda_fa_4_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_58_0/A dadda_fa_5_57_1/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$310 final_adder.U$$312/B final_adder.U$$310/B VGND VGND VPWR VPWR
+ final_adder.U$$436/B sky130_fd_sc_hd__and2_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$321 final_adder.U$$320/B final_adder.U$$195/X final_adder.U$$193/X
+ VGND VGND VPWR VPWR final_adder.U$$321/X sky130_fd_sc_hd__a21o_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$332 final_adder.U$$334/B final_adder.U$$332/B VGND VGND VPWR VPWR
+ final_adder.U$$458/B sky130_fd_sc_hd__and2_1
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$343 final_adder.U$$342/B final_adder.U$$217/X final_adder.U$$215/X
+ VGND VGND VPWR VPWR final_adder.U$$343/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$354 final_adder.U$$356/B final_adder.U$$354/B VGND VGND VPWR VPWR
+ final_adder.U$$480/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$365 final_adder.U$$364/B final_adder.U$$239/X final_adder.U$$237/X
+ VGND VGND VPWR VPWR final_adder.U$$365/X sky130_fd_sc_hd__a21o_1
XU$$204 U$$204/A U$$220/B VGND VGND VPWR VPWR U$$204/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$376 final_adder.U$$378/B final_adder.U$$376/B VGND VGND VPWR VPWR
+ final_adder.U$$498/A sky130_fd_sc_hd__and2_1
XU$$215 U$$215/A1 U$$219/A2 U$$215/B1 U$$219/B2 VGND VGND VPWR VPWR U$$216/A sky130_fd_sc_hd__a22o_1
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$387 final_adder.U$$386/B final_adder.U$$265/X final_adder.U$$261/X
+ VGND VGND VPWR VPWR final_adder.U$$387/X sky130_fd_sc_hd__a21o_1
XU$$226 U$$226/A U$$230/B VGND VGND VPWR VPWR U$$226/X sky130_fd_sc_hd__xor2_1
XFILLER_45_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$398 final_adder.U$$402/B final_adder.U$$398/B VGND VGND VPWR VPWR
+ final_adder.U$$522/B sky130_fd_sc_hd__and2_1
XU$$237 U$$922/A1 U$$259/A2 U$$922/B1 U$$259/B2 VGND VGND VPWR VPWR U$$238/A sky130_fd_sc_hd__a22o_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$248 U$$248/A U$$254/B VGND VGND VPWR VPWR U$$248/X sky130_fd_sc_hd__xor2_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$259 U$$944/A1 U$$259/A2 U$$944/B1 U$$259/B2 VGND VGND VPWR VPWR U$$260/A sky130_fd_sc_hd__a22o_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$9 U$$9/A U$$9/B VGND VGND VPWR VPWR U$$9/X sky130_fd_sc_hd__xor2_1
XFILLER_153_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_75_0 U$$821/Y U$$955/X U$$1088/X VGND VGND VPWR VPWR dadda_fa_1_76_8/A
+ dadda_fa_1_75_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$760 U$$760/A U$$764/B VGND VGND VPWR VPWR U$$760/X sky130_fd_sc_hd__xor2_1
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$771 U$$906/B1 U$$771/A2 U$$773/A1 U$$771/B2 VGND VGND VPWR VPWR U$$772/A sky130_fd_sc_hd__a22o_1
XU$$782 U$$782/A U$$820/B VGND VGND VPWR VPWR U$$782/X sky130_fd_sc_hd__xor2_1
XU$$793 U$$930/A1 U$$809/A2 U$$932/A1 U$$809/B2 VGND VGND VPWR VPWR U$$794/A sky130_fd_sc_hd__a22o_1
XFILLER_91_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_81_1 dadda_fa_5_81_1/A dadda_fa_5_81_1/B dadda_fa_5_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_82_0/B dadda_fa_7_81_0/A sky130_fd_sc_hd__fa_2
XFILLER_145_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_97_1 U$$2728/X U$$2861/X U$$2994/X VGND VGND VPWR VPWR dadda_fa_3_98_0/CIN
+ dadda_fa_3_97_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_74_0 dadda_fa_5_74_0/A dadda_fa_5_74_0/B dadda_fa_5_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_75_0/A dadda_fa_6_74_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_126_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout506 U$$3257/A2 VGND VGND VPWR VPWR U$$3255/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout517 U$$3118/A2 VGND VGND VPWR VPWR U$$3148/A2 sky130_fd_sc_hd__buf_4
Xfanout528 U$$278/X VGND VGND VPWR VPWR U$$362/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_73_8 dadda_fa_1_73_8/A dadda_fa_1_73_8/B dadda_fa_1_73_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_74_3/A dadda_fa_3_73_0/A sky130_fd_sc_hd__fa_2
XFILLER_112_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout539 U$$2844/A2 VGND VGND VPWR VPWR U$$2840/A2 sky130_fd_sc_hd__buf_4
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_66_7 dadda_fa_1_66_7/A dadda_fa_1_66_7/B dadda_fa_1_66_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_67_2/CIN dadda_fa_2_66_5/CIN sky130_fd_sc_hd__fa_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_59_6 U$$3982/X input211/X dadda_fa_1_59_6/CIN VGND VGND VPWR VPWR dadda_fa_2_60_2/B
+ dadda_fa_2_59_5/B sky130_fd_sc_hd__fa_1
XFILLER_67_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_89_0 dadda_fa_7_89_0/A dadda_fa_7_89_0/B dadda_fa_7_89_0/CIN VGND VGND
+ VPWR VPWR _386_/D _257_/D sky130_fd_sc_hd__fa_1
XFILLER_163_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_92_0 dadda_fa_1_92_0/A U$$2053/X U$$2186/X VGND VGND VPWR VPWR dadda_fa_2_93_4/CIN
+ dadda_fa_2_92_5/B sky130_fd_sc_hd__fa_1
XFILLER_150_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4508 U$$4508/A1 U$$4388/X U$$4508/B1 U$$4508/B2 VGND VGND VPWR VPWR U$$4509/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$140 final_adder.U$$140/A final_adder.U$$140/B VGND VGND VPWR VPWR
+ final_adder.U$$268/B sky130_fd_sc_hd__and2_1
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3807 U$$4492/A1 U$$3825/A2 U$$4492/B1 U$$3825/B2 VGND VGND VPWR VPWR U$$3808/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3818 U$$3818/A U$$3828/B VGND VGND VPWR VPWR U$$3818/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$151 final_adder.U$$150/B final_adder.U$$921/B1 final_adder.U$$151/B1
+ VGND VGND VPWR VPWR final_adder.U$$151/X sky130_fd_sc_hd__a21o_1
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3829 U$$4375/B1 U$$3829/A2 U$$4240/B1 U$$3829/B2 VGND VGND VPWR VPWR U$$3830/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$162 final_adder.U$$162/A final_adder.U$$162/B VGND VGND VPWR VPWR
+ final_adder.U$$290/B sky130_fd_sc_hd__and2_1
Xdadda_fa_6_104_0 dadda_fa_6_104_0/A dadda_fa_6_104_0/B dadda_fa_6_104_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_105_0/B dadda_fa_7_104_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$173 final_adder.U$$172/B final_adder.U$$943/B1 final_adder.U$$173/B1
+ VGND VGND VPWR VPWR final_adder.U$$173/X sky130_fd_sc_hd__a21o_1
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$184 final_adder.U$$184/A final_adder.U$$184/B VGND VGND VPWR VPWR
+ final_adder.U$$312/B sky130_fd_sc_hd__and2_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$195 final_adder.U$$194/B final_adder.U$$965/B1 final_adder.U$$195/B1
+ VGND VGND VPWR VPWR final_adder.U$$195/X sky130_fd_sc_hd__a21o_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_24_3 input173/X dadda_fa_3_24_3/B dadda_fa_3_24_3/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_25_1/B dadda_fa_4_24_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_385_ _386_/CLK _385_/D VGND VGND VPWR VPWR _385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_91_0 dadda_fa_6_91_0/A dadda_fa_6_91_0/B dadda_fa_6_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_92_0/B dadda_fa_7_91_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_154_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_69_5 dadda_fa_2_69_5/A dadda_fa_2_69_5/B dadda_fa_2_69_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_2/A dadda_fa_4_69_0/A sky130_fd_sc_hd__fa_1
XFILLER_1_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput180 c[30] VGND VGND VPWR VPWR input180/X sky130_fd_sc_hd__clkbuf_2
Xinput191 c[40] VGND VGND VPWR VPWR input191/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$590 U$$864/A1 U$$630/A2 U$$864/B1 U$$630/B2 VGND VGND VPWR VPWR U$$591/A sky130_fd_sc_hd__a22o_1
XFILLER_108_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_71_5 U$$4139/X U$$4272/X U$$4405/X VGND VGND VPWR VPWR dadda_fa_2_72_2/A
+ dadda_fa_2_71_5/A sky130_fd_sc_hd__fa_1
XFILLER_59_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_4 U$$4125/X U$$4258/X U$$4391/X VGND VGND VPWR VPWR dadda_fa_2_65_1/CIN
+ dadda_fa_2_64_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_57_3 U$$2382/X U$$2515/X U$$2648/X VGND VGND VPWR VPWR dadda_fa_2_58_1/B
+ dadda_fa_2_57_4/B sky130_fd_sc_hd__fa_1
XFILLER_27_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_34_2 dadda_fa_4_34_2/A dadda_fa_4_34_2/B dadda_fa_4_34_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_35_0/CIN dadda_fa_5_34_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_957 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_27_1 dadda_fa_4_27_1/A dadda_fa_4_27_1/B dadda_fa_4_27_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_28_0/B dadda_fa_5_27_1/B sky130_fd_sc_hd__fa_1
XFILLER_15_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_170_ _319_/CLK _170_/D VGND VGND VPWR VPWR _170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4305 U$$4440/B1 U$$4381/A2 U$$4307/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4306/A
+ sky130_fd_sc_hd__a22o_1
Xfanout870 U$$1649/X VGND VGND VPWR VPWR U$$1760/B2 sky130_fd_sc_hd__buf_6
XU$$4316 U$$4316/A U$$4368/B VGND VGND VPWR VPWR U$$4316/X sky130_fd_sc_hd__xor2_1
Xfanout881 U$$259/B2 VGND VGND VPWR VPWR U$$219/B2 sky130_fd_sc_hd__buf_4
XU$$4327 U$$4464/A1 U$$4349/A2 U$$4464/B1 U$$4349/B2 VGND VGND VPWR VPWR U$$4328/A
+ sky130_fd_sc_hd__a22o_1
Xfanout892 U$$1480/B2 VGND VGND VPWR VPWR U$$1452/B2 sky130_fd_sc_hd__buf_6
XFILLER_93_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4338 U$$4338/A U$$4360/B VGND VGND VPWR VPWR U$$4338/X sky130_fd_sc_hd__xor2_1
XU$$3604 U$$4426/A1 U$$3604/A2 U$$4428/A1 U$$3604/B2 VGND VGND VPWR VPWR U$$3605/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4349 U$$4349/A1 U$$4349/A2 U$$4349/B1 U$$4349/B2 VGND VGND VPWR VPWR U$$4350/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_3_16_1 U$$438/X U$$571/X VGND VGND VPWR VPWR dadda_fa_4_17_2/A dadda_ha_3_16_1/SUM
+ sky130_fd_sc_hd__ha_1
XU$$3615 U$$3615/A U$$3615/B VGND VGND VPWR VPWR U$$3615/X sky130_fd_sc_hd__xor2_1
XU$$3626 U$$3763/A1 U$$3640/A2 U$$3628/A1 U$$3640/B2 VGND VGND VPWR VPWR U$$3627/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3637 U$$3637/A U$$3641/B VGND VGND VPWR VPWR U$$3637/X sky130_fd_sc_hd__xor2_1
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3648 U$$4470/A1 U$$3696/A2 U$$3650/A1 U$$3696/B2 VGND VGND VPWR VPWR U$$3649/A
+ sky130_fd_sc_hd__a22o_1
XU$$2903 U$$3314/A1 U$$2991/A2 U$$28/A1 U$$2991/B2 VGND VGND VPWR VPWR U$$2904/A sky130_fd_sc_hd__a22o_1
XU$$3659 U$$3659/A U$$3659/B VGND VGND VPWR VPWR U$$3659/X sky130_fd_sc_hd__xor2_1
XU$$2914 U$$2914/A U$$2944/B VGND VGND VPWR VPWR U$$2914/X sky130_fd_sc_hd__xor2_1
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2925 U$$2925/A1 U$$2929/A2 U$$3338/A1 U$$2929/B2 VGND VGND VPWR VPWR U$$2926/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2936 U$$2936/A U$$2938/B VGND VGND VPWR VPWR U$$2936/X sky130_fd_sc_hd__xor2_1
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_22_0 U$$317/X U$$450/X U$$583/X VGND VGND VPWR VPWR dadda_fa_4_23_0/B
+ dadda_fa_4_22_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2947 U$$479/B1 U$$2991/A2 U$$346/A1 U$$2991/B2 VGND VGND VPWR VPWR U$$2948/A sky130_fd_sc_hd__a22o_1
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2958 U$$2958/A U$$3014/A VGND VGND VPWR VPWR U$$2958/X sky130_fd_sc_hd__xor2_1
XU$$2969 U$$3106/A1 U$$2979/A2 U$$3106/B1 U$$2979/B2 VGND VGND VPWR VPWR U$$2970/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_368_ _368_/CLK _368_/D VGND VGND VPWR VPWR _368_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_147_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_299_ _319_/CLK _299_/D VGND VGND VPWR VPWR _299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_81_4 dadda_fa_2_81_4/A dadda_fa_2_81_4/B dadda_fa_2_81_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_1/CIN dadda_fa_3_81_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_74_3 dadda_fa_2_74_3/A dadda_fa_2_74_3/B dadda_fa_2_74_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_1/B dadda_fa_3_74_3/B sky130_fd_sc_hd__fa_1
XFILLER_96_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_67_2 dadda_fa_2_67_2/A dadda_fa_2_67_2/B dadda_fa_2_67_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_1/A dadda_fa_3_67_3/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$909 final_adder.U$$138/A final_adder.U$$847/X final_adder.U$$909/B1
+ VGND VGND VPWR VPWR final_adder.U$$909/X sky130_fd_sc_hd__a21o_1
XFILLER_69_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_44_1 dadda_fa_5_44_1/A dadda_fa_5_44_1/B dadda_fa_5_44_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_45_0/B dadda_fa_7_44_0/A sky130_fd_sc_hd__fa_1
XFILLER_3_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_37_0 dadda_fa_5_37_0/A dadda_fa_5_37_0/B dadda_fa_5_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_38_0/A dadda_fa_6_37_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_25_916 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_111_0 dadda_fa_5_111_0/A dadda_fa_5_111_0/B dadda_fa_5_111_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_112_0/A dadda_fa_6_111_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_146_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$965_1916 VGND VGND VPWR VPWR U$$965_1916/HI U$$965/A1 sky130_fd_sc_hd__conb_1
Xfanout1109 input80/X VGND VGND VPWR VPWR U$$3751/B1 sky130_fd_sc_hd__buf_4
XFILLER_59_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_62_1 U$$2791/X U$$2924/X U$$3057/X VGND VGND VPWR VPWR dadda_fa_2_63_0/CIN
+ dadda_fa_2_62_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_55_0 U$$782/X U$$915/X U$$1048/X VGND VGND VPWR VPWR dadda_fa_2_56_0/B
+ dadda_fa_2_55_3/B sky130_fd_sc_hd__fa_1
XFILLER_74_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1509 U$$1644/A VGND VGND VPWR VPWR U$$1509/Y sky130_fd_sc_hd__inv_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_222_ _353_/CLK _222_/D VGND VGND VPWR VPWR _222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_91_3 dadda_fa_3_91_3/A dadda_fa_3_91_3/B dadda_fa_3_91_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_1/B dadda_fa_4_91_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_84_2 dadda_fa_3_84_2/A dadda_fa_3_84_2/B dadda_fa_3_84_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_1/A dadda_fa_4_84_2/B sky130_fd_sc_hd__fa_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_864 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_77_1 dadda_fa_3_77_1/A dadda_fa_3_77_1/B dadda_fa_3_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_0/CIN dadda_fa_4_77_2/A sky130_fd_sc_hd__fa_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_54_0 dadda_fa_6_54_0/A dadda_fa_6_54_0/B dadda_fa_6_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_55_0/B dadda_fa_7_54_0/CIN sky130_fd_sc_hd__fa_1
Xfanout1610 U$$2175/B1 VGND VGND VPWR VPWR U$$805/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout1621 input116/X VGND VGND VPWR VPWR U$$2312/A1 sky130_fd_sc_hd__buf_2
XFILLER_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1632 U$$4502/A1 VGND VGND VPWR VPWR U$$4365/A1 sky130_fd_sc_hd__buf_4
Xfanout1643 U$$4500/A1 VGND VGND VPWR VPWR U$$3815/A1 sky130_fd_sc_hd__buf_4
Xfanout1654 input113/X VGND VGND VPWR VPWR U$$2578/B1 sky130_fd_sc_hd__buf_8
XU$$4102 U$$4102/A U$$4108/B VGND VGND VPWR VPWR U$$4102/X sky130_fd_sc_hd__xor2_1
Xfanout1665 U$$2711/B1 VGND VGND VPWR VPWR U$$2576/A1 sky130_fd_sc_hd__buf_6
XU$$4113 U$$4247/A U$$4113/B VGND VGND VPWR VPWR U$$4113/X sky130_fd_sc_hd__and2_1
XFILLER_144_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4124 U$$4259/B1 U$$4158/A2 U$$4400/A1 U$$4158/B2 VGND VGND VPWR VPWR U$$4125/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1676 fanout1680/X VGND VGND VPWR VPWR U$$517/B1 sky130_fd_sc_hd__clkbuf_4
XU$$4135 U$$4135/A U$$4159/B VGND VGND VPWR VPWR U$$4135/X sky130_fd_sc_hd__xor2_1
Xfanout1687 U$$1360/B VGND VGND VPWR VPWR U$$1320/B sky130_fd_sc_hd__buf_6
XU$$3401 U$$3401/A U$$3417/B VGND VGND VPWR VPWR U$$3401/X sky130_fd_sc_hd__xor2_1
XU$$4146 U$$4283/A1 U$$4190/A2 U$$4422/A1 U$$4190/B2 VGND VGND VPWR VPWR U$$4147/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1698 U$$3713/B1 VGND VGND VPWR VPWR U$$562/B1 sky130_fd_sc_hd__buf_2
XU$$4157 U$$4157/A U$$4175/B VGND VGND VPWR VPWR U$$4157/X sky130_fd_sc_hd__xor2_1
XU$$3412 U$$3684/B1 U$$3416/A2 U$$3551/A1 U$$3416/B2 VGND VGND VPWR VPWR U$$3413/A
+ sky130_fd_sc_hd__a22o_1
XU$$4168 U$$4440/B1 U$$4174/A2 U$$4307/A1 U$$4174/B2 VGND VGND VPWR VPWR U$$4169/A
+ sky130_fd_sc_hd__a22o_1
XU$$3423 U$$3423/A U$$3424/A VGND VGND VPWR VPWR U$$3423/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_113_2 dadda_fa_4_113_2/A dadda_fa_4_113_2/B dadda_fa_4_113_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_114_0/CIN dadda_fa_5_113_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_168_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3434 U$$3434/A U$$3468/B VGND VGND VPWR VPWR U$$3434/X sky130_fd_sc_hd__xor2_1
XFILLER_93_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4179 U$$4179/A U$$4231/B VGND VGND VPWR VPWR U$$4179/X sky130_fd_sc_hd__xor2_1
XU$$2700 U$$2700/A U$$2708/B VGND VGND VPWR VPWR U$$2700/X sky130_fd_sc_hd__xor2_1
XU$$3445 U$$3580/B1 U$$3523/A2 U$$4406/A1 U$$3523/B2 VGND VGND VPWR VPWR U$$3446/A
+ sky130_fd_sc_hd__a22o_1
XU$$3456 U$$3456/A U$$3468/B VGND VGND VPWR VPWR U$$3456/X sky130_fd_sc_hd__xor2_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2711 U$$2711/A1 U$$2711/A2 U$$2711/B1 U$$2711/B2 VGND VGND VPWR VPWR U$$2712/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3467 U$$4426/A1 U$$3471/A2 U$$4428/A1 U$$3471/B2 VGND VGND VPWR VPWR U$$3468/A
+ sky130_fd_sc_hd__a22o_1
XU$$2722 U$$2722/A U$$2738/B VGND VGND VPWR VPWR U$$2722/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_106_1 dadda_fa_4_106_1/A dadda_fa_4_106_1/B dadda_fa_4_106_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_107_0/B dadda_fa_5_106_1/B sky130_fd_sc_hd__fa_1
XU$$2733 U$$3418/A1 U$$2733/A2 U$$3418/B1 U$$2733/B2 VGND VGND VPWR VPWR U$$2734/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3478 U$$3478/A U$$3482/B VGND VGND VPWR VPWR U$$3478/X sky130_fd_sc_hd__xor2_1
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2744 U$$2742/Y input35/X U$$2745/A2 U$$2743/X U$$2740/Y VGND VGND VPWR VPWR U$$2744/X
+ sky130_fd_sc_hd__a32o_2
XU$$3489 U$$3763/A1 U$$3505/A2 U$$3628/A1 U$$3505/B2 VGND VGND VPWR VPWR U$$3490/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2755 U$$2755/A U$$2799/B VGND VGND VPWR VPWR U$$2755/X sky130_fd_sc_hd__xor2_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2766 U$$709/B1 U$$2856/A2 U$$576/A1 U$$2856/B2 VGND VGND VPWR VPWR U$$2767/A sky130_fd_sc_hd__a22o_1
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2777 U$$2777/A U$$2811/B VGND VGND VPWR VPWR U$$2777/X sky130_fd_sc_hd__xor2_1
XU$$2788 U$$2925/A1 U$$2804/A2 U$$3338/A1 U$$2804/B2 VGND VGND VPWR VPWR U$$2789/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2799 U$$2799/A U$$2799/B VGND VGND VPWR VPWR U$$2799/X sky130_fd_sc_hd__xor2_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_127_0 dadda_fa_7_127_0/A dadda_fa_7_127_0/B dadda_fa_7_127_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_127_0/COUT _295_/D sky130_fd_sc_hd__fa_1
XFILLER_105_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_72_0 dadda_fa_2_72_0/A dadda_fa_2_72_0/B dadda_fa_2_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_0/B dadda_fa_3_72_2/B sky130_fd_sc_hd__fa_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$706 final_adder.U$$706/A final_adder.U$$706/B VGND VGND VPWR VPWR
+ final_adder.U$$786/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$717 final_adder.U$$716/B final_adder.U$$613/X final_adder.U$$597/X
+ VGND VGND VPWR VPWR final_adder.U$$717/X sky130_fd_sc_hd__a21o_1
XFILLER_84_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3990 U$$3990/A U$$4026/B VGND VGND VPWR VPWR U$$3990/X sky130_fd_sc_hd__xor2_1
XFILLER_80_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_94_1 dadda_fa_4_94_1/A dadda_fa_4_94_1/B dadda_fa_4_94_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_95_0/B dadda_fa_5_94_1/B sky130_fd_sc_hd__fa_1
XFILLER_106_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_71_0 dadda_fa_7_71_0/A dadda_fa_7_71_0/B dadda_fa_7_71_0/CIN VGND VGND
+ VPWR VPWR _368_/D _239_/D sky130_fd_sc_hd__fa_1
XFILLER_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_87_0 dadda_fa_4_87_0/A dadda_fa_4_87_0/B dadda_fa_4_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_88_0/A dadda_fa_5_87_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_108_3 U$$4479/X input138/X dadda_fa_3_108_3/CIN VGND VGND VPWR VPWR dadda_fa_4_109_1/B
+ dadda_fa_4_108_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput270 output270/A VGND VGND VPWR VPWR o[111] sky130_fd_sc_hd__buf_2
Xoutput281 output281/A VGND VGND VPWR VPWR o[121] sky130_fd_sc_hd__buf_2
Xoutput292 output292/A VGND VGND VPWR VPWR o[16] sky130_fd_sc_hd__buf_2
XFILLER_88_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2007 U$$2007/A U$$2007/B VGND VGND VPWR VPWR U$$2007/X sky130_fd_sc_hd__xor2_1
XFILLER_16_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2018 U$$3249/B1 U$$2052/A2 U$$4486/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2019/A
+ sky130_fd_sc_hd__a22o_1
XU$$2029 U$$2029/A U$$2043/B VGND VGND VPWR VPWR U$$2029/X sky130_fd_sc_hd__xor2_1
XFILLER_28_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1306 U$$1306/A U$$1320/B VGND VGND VPWR VPWR U$$1306/X sky130_fd_sc_hd__xor2_1
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1317 U$$3920/A1 U$$1353/A2 U$$906/B1 U$$1353/B2 VGND VGND VPWR VPWR U$$1318/A
+ sky130_fd_sc_hd__a22o_1
XU$$1328 U$$1328/A U$$1328/B VGND VGND VPWR VPWR U$$1328/X sky130_fd_sc_hd__xor2_1
XU$$1339 U$$2707/B1 U$$1367/A2 U$$2574/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1340/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_924 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_205_ _344_/CLK _205_/D VGND VGND VPWR VPWR _205_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$1100 final_adder.U$$178/A final_adder.U$$887/X VGND VGND VPWR VPWR
+ output358/A sky130_fd_sc_hd__xor2_1
XFILLER_128_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1111 final_adder.U$$168/B final_adder.U$$939/X VGND VGND VPWR VPWR
+ output370/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1122 final_adder.U$$156/A final_adder.U$$865/X VGND VGND VPWR VPWR
+ output382/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1133 final_adder.U$$146/B final_adder.U$$917/X VGND VGND VPWR VPWR
+ output267/A sky130_fd_sc_hd__xor2_1
XFILLER_8_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1144 final_adder.U$$134/A final_adder.U$$843/X VGND VGND VPWR VPWR
+ output280/A sky130_fd_sc_hd__xor2_1
XFILLER_116_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1440 U$$2273/B VGND VGND VPWR VPWR U$$2269/B sky130_fd_sc_hd__buf_8
XFILLER_78_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1451 U$$2148/B VGND VGND VPWR VPWR U$$2106/B sky130_fd_sc_hd__buf_6
XFILLER_93_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1462 U$$2054/A VGND VGND VPWR VPWR U$$2015/B sky130_fd_sc_hd__buf_6
Xfanout1473 U$$1874/B VGND VGND VPWR VPWR U$$1910/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_51_5 dadda_fa_2_51_5/A dadda_fa_2_51_5/B dadda_fa_2_51_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_2/A dadda_fa_4_51_0/A sky130_fd_sc_hd__fa_2
Xfanout1484 U$$1781/A VGND VGND VPWR VPWR U$$1761/B sky130_fd_sc_hd__buf_6
XFILLER_94_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1495 input16/X VGND VGND VPWR VPWR U$$1626/B sky130_fd_sc_hd__buf_8
XFILLER_54_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_44_4 dadda_fa_2_44_4/A dadda_fa_2_44_4/B dadda_fa_2_44_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_45_1/CIN dadda_fa_3_44_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3220 U$$3220/A U$$3287/A VGND VGND VPWR VPWR U$$3220/X sky130_fd_sc_hd__xor2_1
XU$$3231 U$$3503/B1 U$$3241/A2 U$$3370/A1 U$$3241/B2 VGND VGND VPWR VPWR U$$3232/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_6_3_0 U$$13/X U$$146/X VGND VGND VPWR VPWR dadda_fa_7_4_0/B dadda_ha_6_3_0/SUM
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$13 _309_/Q _181_/Q VGND VGND VPWR VPWR final_adder.U$$243/B1 final_adder.U$$242/B
+ sky130_fd_sc_hd__ha_1
XU$$3242 U$$3242/A U$$3242/B VGND VGND VPWR VPWR U$$3242/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$24 _320_/Q _192_/Q VGND VGND VPWR VPWR final_adder.U$$231/A2 final_adder.U$$230/A
+ sky130_fd_sc_hd__ha_1
XU$$3253 U$$4349/A1 U$$3283/A2 U$$4349/B1 U$$3283/B2 VGND VGND VPWR VPWR U$$3254/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$35 _331_/Q _203_/Q VGND VGND VPWR VPWR final_adder.U$$221/B1 final_adder.U$$220/B
+ sky130_fd_sc_hd__ha_1
XU$$3264 U$$3264/A U$$3284/B VGND VGND VPWR VPWR U$$3264/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_37_3 U$$1943/X U$$2076/X U$$2209/X VGND VGND VPWR VPWR dadda_fa_3_38_1/B
+ dadda_fa_3_37_3/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$46 _342_/Q _214_/Q VGND VGND VPWR VPWR final_adder.U$$979/B1 final_adder.U$$208/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$57 _353_/Q _225_/Q VGND VGND VPWR VPWR final_adder.U$$199/B1 final_adder.U$$198/B
+ sky130_fd_sc_hd__ha_1
XU$$2530 U$$3763/A1 U$$2574/A2 U$$3628/A1 U$$2574/B2 VGND VGND VPWR VPWR U$$2531/A
+ sky130_fd_sc_hd__a22o_1
XU$$3275 U$$3960/A1 U$$3285/A2 U$$3960/B1 U$$3285/B2 VGND VGND VPWR VPWR U$$3276/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2541 U$$2541/A U$$2541/B VGND VGND VPWR VPWR U$$2541/X sky130_fd_sc_hd__xor2_1
XU$$3286 U$$3286/A U$$3286/B VGND VGND VPWR VPWR U$$3286/X sky130_fd_sc_hd__xor2_1
XU$$3297 U$$3297/A U$$3335/B VGND VGND VPWR VPWR U$$3297/X sky130_fd_sc_hd__xor2_1
XU$$2552 U$$4196/A1 U$$2598/A2 U$$4196/B1 U$$2598/B2 VGND VGND VPWR VPWR U$$2553/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$68 _364_/Q _236_/Q VGND VGND VPWR VPWR final_adder.U$$957/B1 final_adder.U$$186/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$79 _375_/Q _247_/Q VGND VGND VPWR VPWR final_adder.U$$177/B1 final_adder.U$$176/B
+ sky130_fd_sc_hd__ha_1
XU$$2563 U$$2563/A U$$2575/B VGND VGND VPWR VPWR U$$2563/X sky130_fd_sc_hd__xor2_1
XU$$2574 U$$2574/A1 U$$2574/A2 U$$2576/A1 U$$2574/B2 VGND VGND VPWR VPWR U$$2575/A
+ sky130_fd_sc_hd__a22o_1
XU$$1840 U$$1840/A U$$1854/B VGND VGND VPWR VPWR U$$1840/X sky130_fd_sc_hd__xor2_1
XU$$2585 U$$2585/A U$$2591/B VGND VGND VPWR VPWR U$$2585/X sky130_fd_sc_hd__xor2_1
XU$$1851 U$$479/B1 U$$1881/A2 U$$346/A1 U$$1881/B2 VGND VGND VPWR VPWR U$$1852/A sky130_fd_sc_hd__a22o_1
XU$$2596 U$$3418/A1 U$$2600/A2 U$$954/A1 U$$2600/B2 VGND VGND VPWR VPWR U$$2597/A
+ sky130_fd_sc_hd__a22o_1
XU$$1862 U$$1862/A U$$1874/B VGND VGND VPWR VPWR U$$1862/X sky130_fd_sc_hd__xor2_1
XU$$1873 U$$503/A1 U$$1909/A2 U$$505/A1 U$$1909/B2 VGND VGND VPWR VPWR U$$1874/A sky130_fd_sc_hd__a22o_1
XU$$1884 U$$1884/A U$$1916/B VGND VGND VPWR VPWR U$$1884/X sky130_fd_sc_hd__xor2_1
XU$$1895 U$$388/A1 U$$1909/A2 U$$2443/B1 U$$1909/B2 VGND VGND VPWR VPWR U$$1896/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_957 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$503 final_adder.U$$498/A final_adder.U$$381/X final_adder.U$$377/X
+ VGND VGND VPWR VPWR final_adder.U$$503/X sky130_fd_sc_hd__a21o_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$514 final_adder.U$$522/B final_adder.U$$514/B VGND VGND VPWR VPWR
+ final_adder.U$$634/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$525 final_adder.U$$524/B final_adder.U$$409/X final_adder.U$$401/X
+ VGND VGND VPWR VPWR final_adder.U$$525/X sky130_fd_sc_hd__a21o_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$536 final_adder.U$$544/B final_adder.U$$536/B VGND VGND VPWR VPWR
+ final_adder.U$$656/B sky130_fd_sc_hd__and2_1
XFILLER_96_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$547 final_adder.U$$546/B final_adder.U$$431/X final_adder.U$$423/X
+ VGND VGND VPWR VPWR final_adder.U$$547/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$558 final_adder.U$$566/B final_adder.U$$558/B VGND VGND VPWR VPWR
+ final_adder.U$$678/B sky130_fd_sc_hd__and2_1
XFILLER_45_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$569 final_adder.U$$568/B final_adder.U$$453/X final_adder.U$$445/X
+ VGND VGND VPWR VPWR final_adder.U$$569/X sky130_fd_sc_hd__a21o_1
XU$$408 U$$545/A1 U$$408/A2 U$$408/B1 U$$408/B2 VGND VGND VPWR VPWR U$$409/A sky130_fd_sc_hd__a22o_1
XFILLER_72_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$419 U$$965/B1 U$$447/A2 U$$10/A1 U$$447/B2 VGND VGND VPWR VPWR U$$420/A sky130_fd_sc_hd__a22o_1
XFILLER_38_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_113_1 U$$3824/X U$$3957/X U$$4090/X VGND VGND VPWR VPWR dadda_fa_4_114_2/A
+ dadda_fa_4_113_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_147_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_106_0 U$$3544/X U$$3677/X U$$3810/X VGND VGND VPWR VPWR dadda_fa_4_107_0/B
+ dadda_fa_4_106_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_54_3 dadda_fa_3_54_3/A dadda_fa_3_54_3/B dadda_fa_3_54_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_1/B dadda_fa_4_54_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_47_2 dadda_fa_3_47_2/A dadda_fa_3_47_2/B dadda_fa_3_47_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_1/A dadda_fa_4_47_2/B sky130_fd_sc_hd__fa_1
XFILLER_48_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$920 U$$920/A1 U$$956/A2 U$$920/B1 U$$956/B2 VGND VGND VPWR VPWR U$$921/A sky130_fd_sc_hd__a22o_1
XFILLER_16_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$931 U$$931/A U$$959/A VGND VGND VPWR VPWR U$$931/X sky130_fd_sc_hd__xor2_1
XFILLER_28_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$942 U$$942/A1 U$$942/A2 U$$944/A1 U$$942/B2 VGND VGND VPWR VPWR U$$943/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_17_0 dadda_fa_6_17_0/A dadda_fa_6_17_0/B dadda_fa_6_17_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_18_0/B dadda_fa_7_17_0/CIN sky130_fd_sc_hd__fa_1
XU$$953 U$$953/A U$$955/B VGND VGND VPWR VPWR U$$953/X sky130_fd_sc_hd__xor2_1
XU$$964 U$$962/B U$$943/B input6/X U$$959/Y VGND VGND VPWR VPWR U$$964/X sky130_fd_sc_hd__a22o_4
XU$$1103 U$$1103/A U$$1171/B VGND VGND VPWR VPWR U$$1103/X sky130_fd_sc_hd__xor2_1
XU$$1114 U$$3030/B1 U$$1170/A2 U$$2897/A1 U$$1170/B2 VGND VGND VPWR VPWR U$$1115/A
+ sky130_fd_sc_hd__a22o_1
XU$$975 U$$975/A1 U$$979/A2 U$$18/A1 U$$979/B2 VGND VGND VPWR VPWR U$$976/A sky130_fd_sc_hd__a22o_1
XU$$1125 U$$1125/A U$$1163/B VGND VGND VPWR VPWR U$$1125/X sky130_fd_sc_hd__xor2_1
XU$$986 U$$986/A U$$990/B VGND VGND VPWR VPWR U$$986/X sky130_fd_sc_hd__xor2_1
XU$$997 U$$997/A1 U$$997/A2 U$$997/B1 U$$997/B2 VGND VGND VPWR VPWR U$$998/A sky130_fd_sc_hd__a22o_1
XU$$1136 U$$314/A1 U$$1174/A2 U$$42/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1137/A sky130_fd_sc_hd__a22o_1
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1147 U$$1147/A U$$1171/B VGND VGND VPWR VPWR U$$1147/X sky130_fd_sc_hd__xor2_1
XU$$1158 U$$62/A1 U$$1164/A2 U$$64/A1 U$$1164/B2 VGND VGND VPWR VPWR U$$1159/A sky130_fd_sc_hd__a22o_1
XU$$1169 U$$1169/A U$$1189/B VGND VGND VPWR VPWR U$$1169/X sky130_fd_sc_hd__xor2_1
XFILLER_129_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1270 U$$4159/B VGND VGND VPWR VPWR U$$4133/B sky130_fd_sc_hd__clkbuf_8
Xfanout1281 input56/X VGND VGND VPWR VPWR U$$353/B sky130_fd_sc_hd__buf_4
Xfanout1292 fanout1299/X VGND VGND VPWR VPWR U$$4040/B sky130_fd_sc_hd__buf_6
XFILLER_82_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_42_1 U$$2352/X U$$2485/X U$$2618/X VGND VGND VPWR VPWR dadda_fa_3_43_0/CIN
+ dadda_fa_3_42_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3050 U$$721/A1 U$$3072/A2 U$$721/B1 U$$3072/B2 VGND VGND VPWR VPWR U$$3051/A sky130_fd_sc_hd__a22o_1
XFILLER_35_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3061 U$$3061/A U$$3061/B VGND VGND VPWR VPWR U$$3061/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_35_0 U$$343/X U$$476/X U$$609/X VGND VGND VPWR VPWR dadda_fa_3_36_0/B
+ dadda_fa_3_35_2/B sky130_fd_sc_hd__fa_1
XU$$3072 U$$3072/A1 U$$3072/A2 U$$3072/B1 U$$3072/B2 VGND VGND VPWR VPWR U$$3073/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3083 U$$3083/A U$$3119/B VGND VGND VPWR VPWR U$$3083/X sky130_fd_sc_hd__xor2_1
XU$$3094 U$$3503/B1 U$$3108/A2 U$$3370/A1 U$$3108/B2 VGND VGND VPWR VPWR U$$3095/A
+ sky130_fd_sc_hd__a22o_1
XU$$2360 U$$2360/A U$$2396/B VGND VGND VPWR VPWR U$$2360/X sky130_fd_sc_hd__xor2_1
XU$$2371 U$$2780/B1 U$$2413/A2 U$$2647/A1 U$$2413/B2 VGND VGND VPWR VPWR U$$2372/A
+ sky130_fd_sc_hd__a22o_1
XU$$2382 U$$2382/A U$$2416/B VGND VGND VPWR VPWR U$$2382/X sky130_fd_sc_hd__xor2_1
XU$$2393 U$$2665/B1 U$$2395/A2 U$$66/A1 U$$2395/B2 VGND VGND VPWR VPWR U$$2394/A sky130_fd_sc_hd__a22o_1
XFILLER_50_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1670 U$$709/B1 U$$1702/A2 U$$576/A1 U$$1702/B2 VGND VGND VPWR VPWR U$$1671/A sky130_fd_sc_hd__a22o_1
XFILLER_22_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1681 U$$1681/A U$$1703/B VGND VGND VPWR VPWR U$$1681/X sky130_fd_sc_hd__xor2_1
XFILLER_167_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1692 U$$596/A1 U$$1696/A2 U$$596/B1 U$$1696/B2 VGND VGND VPWR VPWR U$$1693/A sky130_fd_sc_hd__a22o_1
XFILLER_147_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_87_3 U$$2841/X U$$2974/X U$$3107/X VGND VGND VPWR VPWR dadda_fa_2_88_4/A
+ dadda_fa_2_87_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_116_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_64_2 dadda_fa_4_64_2/A dadda_fa_4_64_2/B dadda_fa_4_64_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_65_0/CIN dadda_fa_5_64_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_162_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_57_1 dadda_fa_4_57_1/A dadda_fa_4_57_1/B dadda_fa_4_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_58_0/B dadda_fa_5_57_1/B sky130_fd_sc_hd__fa_1
XFILLER_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$300 final_adder.U$$302/B final_adder.U$$300/B VGND VGND VPWR VPWR
+ final_adder.U$$426/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$311 final_adder.U$$310/B final_adder.U$$185/X final_adder.U$$183/X
+ VGND VGND VPWR VPWR final_adder.U$$311/X sky130_fd_sc_hd__a21o_1
XFILLER_97_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_34_0 dadda_fa_7_34_0/A dadda_fa_7_34_0/B dadda_fa_7_34_0/CIN VGND VGND
+ VPWR VPWR _331_/D _202_/D sky130_fd_sc_hd__fa_2
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$322 final_adder.U$$324/B final_adder.U$$322/B VGND VGND VPWR VPWR
+ final_adder.U$$448/B sky130_fd_sc_hd__and2_1
XFILLER_57_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$333 final_adder.U$$332/B final_adder.U$$207/X final_adder.U$$205/X
+ VGND VGND VPWR VPWR final_adder.U$$333/X sky130_fd_sc_hd__a21o_1
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$344 final_adder.U$$346/B final_adder.U$$344/B VGND VGND VPWR VPWR
+ final_adder.U$$470/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$355 final_adder.U$$354/B final_adder.U$$229/X final_adder.U$$227/X
+ VGND VGND VPWR VPWR final_adder.U$$355/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$366 final_adder.U$$368/B final_adder.U$$366/B VGND VGND VPWR VPWR
+ final_adder.U$$492/B sky130_fd_sc_hd__and2_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$205 U$$616/A1 U$$207/A2 U$$481/A1 U$$207/B2 VGND VGND VPWR VPWR U$$206/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$377 final_adder.U$$376/B final_adder.U$$251/X final_adder.U$$249/X
+ VGND VGND VPWR VPWR final_adder.U$$377/X sky130_fd_sc_hd__a21o_1
XU$$216 U$$216/A U$$220/B VGND VGND VPWR VPWR U$$216/X sky130_fd_sc_hd__xor2_1
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$388 final_adder.U$$392/B final_adder.U$$388/B VGND VGND VPWR VPWR
+ final_adder.U$$512/B sky130_fd_sc_hd__and2_1
XU$$227 U$$90/A1 U$$229/A2 U$$92/A1 U$$229/B2 VGND VGND VPWR VPWR U$$228/A sky130_fd_sc_hd__a22o_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$399 final_adder.U$$398/B final_adder.U$$277/X final_adder.U$$273/X
+ VGND VGND VPWR VPWR final_adder.U$$399/X sky130_fd_sc_hd__a21o_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$238 U$$238/A U$$260/B VGND VGND VPWR VPWR U$$238/X sky130_fd_sc_hd__xor2_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$249 U$$384/B1 U$$253/A2 U$$251/A1 U$$253/B2 VGND VGND VPWR VPWR U$$250/A sky130_fd_sc_hd__a22o_1
XFILLER_26_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_866 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_124_0_1941 VGND VGND VPWR VPWR dadda_fa_5_124_0/A dadda_fa_5_124_0_1941/LO
+ sky130_fd_sc_hd__conb_1
Xdadda_fa_0_75_1 U$$1221/X U$$1354/X U$$1487/X VGND VGND VPWR VPWR dadda_fa_1_76_8/B
+ dadda_fa_2_75_0/A sky130_fd_sc_hd__fa_1
XFILLER_49_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_52_0 dadda_fa_3_52_0/A dadda_fa_3_52_0/B dadda_fa_3_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_0/B dadda_fa_4_52_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_121_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_68_0 dadda_fa_0_68_0/A U$$409/X U$$542/X VGND VGND VPWR VPWR dadda_fa_1_69_5/CIN
+ dadda_fa_1_68_7/B sky130_fd_sc_hd__fa_1
XFILLER_36_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$750 U$$750/A U$$768/B VGND VGND VPWR VPWR U$$750/X sky130_fd_sc_hd__xor2_1
XU$$761 U$$898/A1 U$$763/A2 U$$900/A1 U$$763/B2 VGND VGND VPWR VPWR U$$762/A sky130_fd_sc_hd__a22o_1
XU$$772 U$$772/A U$$774/B VGND VGND VPWR VPWR U$$772/X sky130_fd_sc_hd__xor2_1
XFILLER_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$783 U$$783/A1 U$$817/A2 U$$783/B1 U$$817/B2 VGND VGND VPWR VPWR U$$784/A sky130_fd_sc_hd__a22o_1
XFILLER_50_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$794 U$$794/A U$$804/B VGND VGND VPWR VPWR U$$794/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_97_2 U$$3127/X U$$3260/X U$$3393/X VGND VGND VPWR VPWR dadda_fa_3_98_1/A
+ dadda_fa_3_97_3/A sky130_fd_sc_hd__fa_1
XFILLER_145_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_74_1 dadda_fa_5_74_1/A dadda_fa_5_74_1/B dadda_fa_5_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_75_0/B dadda_fa_7_74_0/A sky130_fd_sc_hd__fa_1
XFILLER_126_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_67_0 dadda_fa_5_67_0/A dadda_fa_5_67_0/B dadda_fa_5_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_68_0/A dadda_fa_6_67_0/CIN sky130_fd_sc_hd__fa_1
Xfanout507 U$$3251/A2 VGND VGND VPWR VPWR U$$3283/A2 sky130_fd_sc_hd__buf_4
Xfanout518 U$$3118/A2 VGND VGND VPWR VPWR U$$3144/A2 sky130_fd_sc_hd__buf_2
Xfanout529 U$$278/X VGND VGND VPWR VPWR U$$352/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_66_8 dadda_fa_1_66_8/A dadda_fa_1_66_8/B dadda_fa_1_66_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_67_3/A dadda_fa_3_66_0/A sky130_fd_sc_hd__fa_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_59_7 dadda_fa_1_59_7/A dadda_fa_1_59_7/B dadda_fa_1_59_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_60_2/CIN dadda_fa_2_59_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_6_0 input223/X dadda_fa_6_6_0/B dadda_fa_6_6_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_7_7_0/B dadda_fa_7_6_0/CIN sky130_fd_sc_hd__fa_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2190 U$$2190/A U$$2191/A VGND VGND VPWR VPWR U$$2190/X sky130_fd_sc_hd__xor2_1
XFILLER_50_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_92_1 U$$2319/X U$$2452/X U$$2585/X VGND VGND VPWR VPWR dadda_fa_2_93_5/A
+ dadda_fa_2_92_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_123_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_85_0 U$$1506/Y U$$1640/X U$$1773/X VGND VGND VPWR VPWR dadda_fa_2_86_2/B
+ dadda_fa_2_85_4/B sky130_fd_sc_hd__fa_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4509 U$$4509/A U$$4509/B VGND VGND VPWR VPWR U$$4509/X sky130_fd_sc_hd__xor2_1
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$130 final_adder.U$$130/A final_adder.U$$130/B VGND VGND VPWR VPWR
+ final_adder.U$$258/B sky130_fd_sc_hd__and2_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3808 U$$3808/A U$$3835/A VGND VGND VPWR VPWR U$$3808/X sky130_fd_sc_hd__xor2_1
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3819 U$$4365/B1 U$$3829/A2 U$$4367/B1 U$$3829/B2 VGND VGND VPWR VPWR U$$3820/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$141 final_adder.U$$140/B final_adder.U$$911/B1 final_adder.U$$141/B1
+ VGND VGND VPWR VPWR final_adder.U$$141/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$152 final_adder.U$$152/A final_adder.U$$152/B VGND VGND VPWR VPWR
+ final_adder.U$$280/B sky130_fd_sc_hd__and2_1
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$163 final_adder.U$$162/B final_adder.U$$933/B1 final_adder.U$$163/B1
+ VGND VGND VPWR VPWR final_adder.U$$163/X sky130_fd_sc_hd__a21o_1
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$174 final_adder.U$$174/A final_adder.U$$174/B VGND VGND VPWR VPWR
+ final_adder.U$$302/B sky130_fd_sc_hd__and2_1
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$185 final_adder.U$$184/B final_adder.U$$955/B1 final_adder.U$$185/B1
+ VGND VGND VPWR VPWR final_adder.U$$185/X sky130_fd_sc_hd__a21o_1
XFILLER_46_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$196 final_adder.U$$196/A final_adder.U$$196/B VGND VGND VPWR VPWR
+ final_adder.U$$324/B sky130_fd_sc_hd__and2_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_5_126_0 dadda_ha_5_126_0/A U$$4382/X VGND VGND VPWR VPWR dadda_fa_7_127_0/A
+ dadda_fa_7_126_0/A sky130_fd_sc_hd__ha_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_384_ _384_/CLK _384_/D VGND VGND VPWR VPWR _384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_84_0 dadda_fa_6_84_0/A dadda_fa_6_84_0/B dadda_fa_6_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_85_0/B dadda_fa_7_84_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_126_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput170 c[21] VGND VGND VPWR VPWR input170/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput181 c[31] VGND VGND VPWR VPWR input181/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput192 c[41] VGND VGND VPWR VPWR input192/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$580 U$$32/A1 U$$610/A2 U$$32/B1 U$$610/B2 VGND VGND VPWR VPWR U$$581/A sky130_fd_sc_hd__a22o_1
XU$$591 U$$591/A U$$631/B VGND VGND VPWR VPWR U$$591/X sky130_fd_sc_hd__xor2_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_43_clk _218_/CLK VGND VGND VPWR VPWR _345_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_71_6 input225/X dadda_fa_1_71_6/B dadda_fa_1_71_6/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_72_2/B dadda_fa_2_71_5/B sky130_fd_sc_hd__fa_1
XFILLER_99_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_5 input217/X dadda_fa_1_64_5/B dadda_fa_1_64_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_65_2/A dadda_fa_2_64_5/A sky130_fd_sc_hd__fa_1
XFILLER_28_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_57_4 U$$2781/X U$$2914/X U$$3047/X VGND VGND VPWR VPWR dadda_fa_2_58_1/CIN
+ dadda_fa_2_57_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_54_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_27_2 dadda_fa_4_27_2/A dadda_fa_4_27_2/B dadda_fa_4_27_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_28_0/CIN dadda_fa_5_27_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_34_clk _388_/CLK VGND VGND VPWR VPWR _366_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout860 U$$1891/B2 VGND VGND VPWR VPWR U$$1915/B2 sky130_fd_sc_hd__buf_6
XU$$4306 U$$4306/A U$$4384/A VGND VGND VPWR VPWR U$$4306/X sky130_fd_sc_hd__xor2_1
Xfanout871 U$$1593/B2 VGND VGND VPWR VPWR U$$1563/B2 sky130_fd_sc_hd__clkbuf_4
XU$$4317 U$$4454/A1 U$$4325/A2 U$$4456/A1 U$$4325/B2 VGND VGND VPWR VPWR U$$4318/A
+ sky130_fd_sc_hd__a22o_1
Xfanout882 U$$259/B2 VGND VGND VPWR VPWR U$$271/B2 sky130_fd_sc_hd__buf_4
Xfanout893 U$$1502/B2 VGND VGND VPWR VPWR U$$1504/B2 sky130_fd_sc_hd__buf_6
XFILLER_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4328 U$$4328/A U$$4360/B VGND VGND VPWR VPWR U$$4328/X sky130_fd_sc_hd__xor2_1
XU$$4339 U$$4474/B1 U$$4359/A2 U$$4341/A1 U$$4359/B2 VGND VGND VPWR VPWR U$$4340/A
+ sky130_fd_sc_hd__a22o_1
XU$$3605 U$$3605/A U$$3607/B VGND VGND VPWR VPWR U$$3605/X sky130_fd_sc_hd__xor2_1
XU$$3616 U$$3751/B1 U$$3696/A2 U$$3618/A1 U$$3696/B2 VGND VGND VPWR VPWR U$$3617/A
+ sky130_fd_sc_hd__a22o_1
XU$$3627 U$$3627/A U$$3641/B VGND VGND VPWR VPWR U$$3627/X sky130_fd_sc_hd__xor2_1
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3638 U$$3775/A1 U$$3640/A2 U$$3638/B1 U$$3640/B2 VGND VGND VPWR VPWR U$$3639/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2904 U$$2904/A U$$2944/B VGND VGND VPWR VPWR U$$2904/X sky130_fd_sc_hd__xor2_1
XFILLER_73_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3649 U$$3649/A U$$3695/B VGND VGND VPWR VPWR U$$3649/X sky130_fd_sc_hd__xor2_1
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2915 U$$38/A1 U$$2991/A2 U$$40/A1 U$$2991/B2 VGND VGND VPWR VPWR U$$2916/A sky130_fd_sc_hd__a22o_1
XU$$2926 U$$2926/A U$$2926/B VGND VGND VPWR VPWR U$$2926/X sky130_fd_sc_hd__xor2_1
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2937 U$$4442/B1 U$$2937/A2 U$$4309/A1 U$$2937/B2 VGND VGND VPWR VPWR U$$2938/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2948 U$$2948/A U$$2990/B VGND VGND VPWR VPWR U$$2948/X sky130_fd_sc_hd__xor2_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2959 U$$3370/A1 U$$2979/A2 U$$3370/B1 U$$2979/B2 VGND VGND VPWR VPWR U$$2960/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_22_1 U$$716/X U$$849/X U$$982/X VGND VGND VPWR VPWR dadda_fa_4_23_0/CIN
+ dadda_fa_4_22_2/A sky130_fd_sc_hd__fa_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_367_ _367_/CLK _367_/D VGND VGND VPWR VPWR _367_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_159_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_298_ _319_/CLK _298_/D VGND VGND VPWR VPWR _298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_81_5 dadda_fa_2_81_5/A dadda_fa_2_81_5/B dadda_fa_2_81_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_2/A dadda_fa_4_81_0/A sky130_fd_sc_hd__fa_2
XFILLER_138_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_74_4 dadda_fa_2_74_4/A dadda_fa_2_74_4/B dadda_fa_2_74_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_1/CIN dadda_fa_3_74_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_67_3 dadda_fa_2_67_3/A dadda_fa_2_67_3/B dadda_fa_2_67_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_1/B dadda_fa_3_67_3/B sky130_fd_sc_hd__fa_1
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_37_1 dadda_fa_5_37_1/A dadda_fa_5_37_1/B dadda_fa_5_37_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_38_0/B dadda_fa_7_37_0/A sky130_fd_sc_hd__fa_1
XFILLER_83_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_928 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_clk _370_/CLK VGND VGND VPWR VPWR _408_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_111_1 dadda_fa_5_111_1/A dadda_fa_5_111_1/B dadda_fa_5_111_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_112_0/B dadda_fa_7_111_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_104_0 dadda_fa_5_104_0/A dadda_fa_5_104_0/B dadda_fa_5_104_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_105_0/A dadda_fa_6_104_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_62_2 U$$3190/X U$$3323/X U$$3456/X VGND VGND VPWR VPWR dadda_fa_2_63_1/A
+ dadda_fa_2_62_4/A sky130_fd_sc_hd__fa_1
XU$$4389_1841 VGND VGND VPWR VPWR U$$4389_1841/HI U$$4389/B1 sky130_fd_sc_hd__conb_1
XFILLER_170_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_55_1 U$$1181/X U$$1314/X U$$1447/X VGND VGND VPWR VPWR dadda_fa_2_56_0/CIN
+ dadda_fa_2_55_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_4_32_0 dadda_fa_4_32_0/A dadda_fa_4_32_0/B dadda_fa_4_32_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_33_0/A dadda_fa_5_32_1/A sky130_fd_sc_hd__fa_1
XFILLER_74_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_48_0 U$$103/X U$$236/X U$$369/X VGND VGND VPWR VPWR dadda_fa_2_49_1/A
+ dadda_fa_2_48_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_221_ _353_/CLK _221_/D VGND VGND VPWR VPWR _221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_84_3 dadda_fa_3_84_3/A dadda_fa_3_84_3/B dadda_fa_3_84_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_1/B dadda_fa_4_84_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_151_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_77_2 dadda_fa_3_77_2/A dadda_fa_3_77_2/B dadda_fa_3_77_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_1/A dadda_fa_4_77_2/B sky130_fd_sc_hd__fa_1
XFILLER_3_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1600 input119/X VGND VGND VPWR VPWR U$$2729/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1611 U$$2175/B1 VGND VGND VPWR VPWR U$$944/A1 sky130_fd_sc_hd__buf_2
Xfanout1622 U$$2860/A1 VGND VGND VPWR VPWR U$$120/A1 sky130_fd_sc_hd__buf_6
Xfanout1633 U$$4502/A1 VGND VGND VPWR VPWR U$$3817/A1 sky130_fd_sc_hd__buf_4
XFILLER_26_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_47_0 dadda_fa_6_47_0/A dadda_fa_6_47_0/B dadda_fa_6_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_48_0/B dadda_fa_7_47_0/CIN sky130_fd_sc_hd__fa_1
Xfanout1644 U$$4500/A1 VGND VGND VPWR VPWR U$$4226/A1 sky130_fd_sc_hd__buf_2
Xfanout1655 U$$2578/A1 VGND VGND VPWR VPWR U$$934/A1 sky130_fd_sc_hd__buf_4
XU$$4103 U$$4375/B1 U$$4105/A2 U$$4240/B1 U$$4105/B2 VGND VGND VPWR VPWR U$$4104/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4114 U$$4112/Y input57/X U$$4110/A U$$4113/X U$$4110/Y VGND VGND VPWR VPWR U$$4114/X
+ sky130_fd_sc_hd__a32o_2
Xfanout1666 U$$4494/A1 VGND VGND VPWR VPWR U$$521/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout1677 fanout1680/X VGND VGND VPWR VPWR U$$4081/A1 sky130_fd_sc_hd__buf_4
XU$$4125 U$$4125/A U$$4133/B VGND VGND VPWR VPWR U$$4125/X sky130_fd_sc_hd__xor2_1
Xfanout1688 U$$1364/B VGND VGND VPWR VPWR U$$1370/A sky130_fd_sc_hd__buf_4
XU$$4136 U$$985/A1 U$$4244/A2 U$$987/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4137/A sky130_fd_sc_hd__a22o_1
Xfanout690 U$$4325/B2 VGND VGND VPWR VPWR U$$4369/B2 sky130_fd_sc_hd__buf_2
XU$$3402 U$$3948/B1 U$$3418/A2 U$$3815/A1 U$$3418/B2 VGND VGND VPWR VPWR U$$3403/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1699 U$$3713/B1 VGND VGND VPWR VPWR U$$973/B1 sky130_fd_sc_hd__buf_4
XU$$4147 U$$4147/A U$$4191/B VGND VGND VPWR VPWR U$$4147/X sky130_fd_sc_hd__xor2_1
XU$$3413 U$$3413/A U$$3417/B VGND VGND VPWR VPWR U$$3413/X sky130_fd_sc_hd__xor2_1
XU$$4158 U$$4158/A1 U$$4158/A2 U$$4295/B1 U$$4158/B2 VGND VGND VPWR VPWR U$$4159/A
+ sky130_fd_sc_hd__a22o_1
XU$$4169 U$$4169/A U$$4175/B VGND VGND VPWR VPWR U$$4169/X sky130_fd_sc_hd__xor2_1
XU$$3424 U$$3424/A VGND VGND VPWR VPWR U$$3424/Y sky130_fd_sc_hd__inv_1
XU$$3435 U$$3435/A1 U$$3439/A2 U$$971/A1 U$$3439/B2 VGND VGND VPWR VPWR U$$3436/A
+ sky130_fd_sc_hd__a22o_1
XU$$2701 U$$2973/B1 U$$2707/A2 U$$2840/A1 U$$2707/B2 VGND VGND VPWR VPWR U$$2702/A
+ sky130_fd_sc_hd__a22o_1
XU$$3446 U$$3446/A U$$3482/B VGND VGND VPWR VPWR U$$3446/X sky130_fd_sc_hd__xor2_1
XU$$3457 U$$854/A1 U$$3471/A2 U$$3870/A1 U$$3471/B2 VGND VGND VPWR VPWR U$$3458/A
+ sky130_fd_sc_hd__a22o_1
XU$$2712 U$$2712/A U$$2740/A VGND VGND VPWR VPWR U$$2712/X sky130_fd_sc_hd__xor2_1
XFILLER_92_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2723 U$$2860/A1 U$$2737/A2 U$$120/B1 U$$2737/B2 VGND VGND VPWR VPWR U$$2724/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_106_2 dadda_fa_4_106_2/A dadda_fa_4_106_2/B dadda_fa_4_106_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_107_0/CIN dadda_fa_5_106_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3468 U$$3468/A U$$3468/B VGND VGND VPWR VPWR U$$3468/X sky130_fd_sc_hd__xor2_1
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2734 U$$2734/A U$$2738/B VGND VGND VPWR VPWR U$$2734/X sky130_fd_sc_hd__xor2_1
XU$$3479 U$$3751/B1 U$$3523/A2 U$$3618/A1 U$$3523/B2 VGND VGND VPWR VPWR U$$3480/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2745 U$$2743/B U$$2745/A2 input35/X U$$2740/Y VGND VGND VPWR VPWR U$$2745/X sky130_fd_sc_hd__a22o_2
XU$$2756 U$$2891/B1 U$$2798/A2 U$$2758/A1 U$$2798/B2 VGND VGND VPWR VPWR U$$2757/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2767 U$$2767/A U$$2811/B VGND VGND VPWR VPWR U$$2767/X sky130_fd_sc_hd__xor2_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2778 U$$4011/A1 U$$2856/A2 U$$2780/A1 U$$2856/B2 VGND VGND VPWR VPWR U$$2779/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2789 U$$2789/A U$$2805/B VGND VGND VPWR VPWR U$$2789/X sky130_fd_sc_hd__xor2_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_419_ _421_/CLK _419_/D VGND VGND VPWR VPWR _419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_clk _201_/CLK VGND VGND VPWR VPWR _344_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_170_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_72_1 dadda_fa_2_72_1/A dadda_fa_2_72_1/B dadda_fa_2_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_0/CIN dadda_fa_3_72_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_65_0 dadda_fa_2_65_0/A dadda_fa_2_65_0/B dadda_fa_2_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_0/B dadda_fa_3_65_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$707 final_adder.U$$706/B final_adder.U$$603/X final_adder.U$$587/X
+ VGND VGND VPWR VPWR final_adder.U$$707/X sky130_fd_sc_hd__a21o_1
XFILLER_111_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$718 final_adder.U$$718/A final_adder.U$$718/B VGND VGND VPWR VPWR
+ final_adder.U$$798/A sky130_fd_sc_hd__and2_1
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$729 final_adder.U$$712/A final_adder.U$$625/X final_adder.U$$609/X
+ VGND VGND VPWR VPWR final_adder.U$$729/X sky130_fd_sc_hd__a21o_2
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3980 U$$3980/A U$$4006/B VGND VGND VPWR VPWR U$$3980/X sky130_fd_sc_hd__xor2_1
XU$$3991 U$$4400/B1 U$$4025/A2 U$$4265/B1 U$$4025/B2 VGND VGND VPWR VPWR U$$3992/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_94_2 dadda_fa_4_94_2/A dadda_fa_4_94_2/B dadda_fa_4_94_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_95_0/CIN dadda_fa_5_94_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_165_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_87_1 dadda_fa_4_87_1/A dadda_fa_4_87_1/B dadda_fa_4_87_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_88_0/B dadda_fa_5_87_1/B sky130_fd_sc_hd__fa_1
XFILLER_173_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_64_0 dadda_fa_7_64_0/A dadda_fa_7_64_0/B dadda_fa_7_64_0/CIN VGND VGND
+ VPWR VPWR _361_/D _232_/D sky130_fd_sc_hd__fa_1
XFILLER_145_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput260 output260/A VGND VGND VPWR VPWR o[102] sky130_fd_sc_hd__buf_2
Xoutput271 output271/A VGND VGND VPWR VPWR o[112] sky130_fd_sc_hd__buf_2
Xoutput282 output282/A VGND VGND VPWR VPWR o[122] sky130_fd_sc_hd__buf_2
Xoutput293 output293/A VGND VGND VPWR VPWR o[17] sky130_fd_sc_hd__buf_2
XFILLER_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2008 U$$88/B1 U$$2022/A2 U$$503/A1 U$$2022/B2 VGND VGND VPWR VPWR U$$2009/A sky130_fd_sc_hd__a22o_1
XFILLER_43_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2019 U$$2019/A U$$2053/B VGND VGND VPWR VPWR U$$2019/X sky130_fd_sc_hd__xor2_1
XU$$1307 U$$74/A1 U$$1309/A2 U$$76/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1308/A sky130_fd_sc_hd__a22o_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1318 U$$1318/A U$$1320/B VGND VGND VPWR VPWR U$$1318/X sky130_fd_sc_hd__xor2_1
XFILLER_71_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1329 U$$96/A1 U$$1367/A2 U$$98/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1330/A sky130_fd_sc_hd__a22o_1
XFILLER_43_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_204_ _344_/CLK _204_/D VGND VGND VPWR VPWR _204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1101 final_adder.U$$178/B final_adder.U$$949/X VGND VGND VPWR VPWR
+ output359/A sky130_fd_sc_hd__xor2_1
XFILLER_12_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1112 final_adder.U$$166/A final_adder.U$$875/X VGND VGND VPWR VPWR
+ output371/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1123 final_adder.U$$156/B final_adder.U$$927/X VGND VGND VPWR VPWR
+ output383/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1134 final_adder.U$$144/A final_adder.U$$853/X VGND VGND VPWR VPWR
+ output269/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1145 final_adder.U$$134/B final_adder.U$$905/X VGND VGND VPWR VPWR
+ output281/A sky130_fd_sc_hd__xor2_1
XFILLER_99_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_82_0 dadda_fa_3_82_0/A dadda_fa_3_82_0/B dadda_fa_3_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_0/B dadda_fa_4_82_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_125_866 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1430 U$$2408/B VGND VGND VPWR VPWR U$$2402/B sky130_fd_sc_hd__buf_6
Xfanout1441 U$$2283/B VGND VGND VPWR VPWR U$$2253/B sky130_fd_sc_hd__buf_6
XFILLER_79_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1452 U$$2140/B VGND VGND VPWR VPWR U$$2148/B sky130_fd_sc_hd__buf_8
Xfanout1463 U$$2031/B VGND VGND VPWR VPWR U$$2043/B sky130_fd_sc_hd__buf_6
Xfanout1474 U$$1874/B VGND VGND VPWR VPWR U$$1918/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1485 input18/X VGND VGND VPWR VPWR U$$1781/A sky130_fd_sc_hd__buf_2
Xfanout1496 U$$1461/B VGND VGND VPWR VPWR U$$1427/B sky130_fd_sc_hd__clkbuf_8
XFILLER_94_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3210 U$$3210/A U$$3210/B VGND VGND VPWR VPWR U$$3210/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_44_5 dadda_fa_2_44_5/A dadda_fa_2_44_5/B dadda_fa_2_44_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_45_2/A dadda_fa_4_44_0/A sky130_fd_sc_hd__fa_1
XU$$3221 U$$3630/B1 U$$3245/A2 U$$3495/B1 U$$3245/B2 VGND VGND VPWR VPWR U$$3222/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_111_0 U$$4485/X input142/X dadda_fa_4_111_0/CIN VGND VGND VPWR VPWR dadda_fa_5_112_0/A
+ dadda_fa_5_111_1/A sky130_fd_sc_hd__fa_1
XFILLER_19_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3232 U$$3232/A U$$3242/B VGND VGND VPWR VPWR U$$3232/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$14 _310_/Q _182_/Q VGND VGND VPWR VPWR final_adder.U$$241/A2 final_adder.U$$240/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$25 _321_/Q _193_/Q VGND VGND VPWR VPWR final_adder.U$$231/B1 final_adder.U$$230/B
+ sky130_fd_sc_hd__ha_1
XU$$3243 U$$3243/A1 U$$3245/A2 U$$3243/B1 U$$3245/B2 VGND VGND VPWR VPWR U$$3244/A
+ sky130_fd_sc_hd__a22o_1
XU$$3254 U$$3254/A U$$3284/B VGND VGND VPWR VPWR U$$3254/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$36 _332_/Q _204_/Q VGND VGND VPWR VPWR final_adder.U$$989/B1 final_adder.U$$218/A
+ sky130_fd_sc_hd__ha_1
XU$$3265 U$$3948/B1 U$$3285/A2 U$$3815/A1 U$$3285/B2 VGND VGND VPWR VPWR U$$3266/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2520 U$$602/A1 U$$2540/A2 U$$3205/B1 U$$2540/B2 VGND VGND VPWR VPWR U$$2521/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_37_4 U$$2342/X U$$2475/X input187/X VGND VGND VPWR VPWR dadda_fa_3_38_1/CIN
+ dadda_fa_3_37_3/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$47 _343_/Q _215_/Q VGND VGND VPWR VPWR final_adder.U$$209/B1 final_adder.U$$208/B
+ sky130_fd_sc_hd__ha_1
XU$$2531 U$$2531/A U$$2575/B VGND VGND VPWR VPWR U$$2531/X sky130_fd_sc_hd__xor2_1
XU$$3276 U$$3276/A U$$3286/B VGND VGND VPWR VPWR U$$3276/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$58 _354_/Q _226_/Q VGND VGND VPWR VPWR final_adder.U$$967/B1 final_adder.U$$196/A
+ sky130_fd_sc_hd__ha_1
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2542 U$$4049/A1 U$$2598/A2 U$$4462/A1 U$$2598/B2 VGND VGND VPWR VPWR U$$2543/A
+ sky130_fd_sc_hd__a22o_1
XU$$3287 U$$3287/A VGND VGND VPWR VPWR U$$3287/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$69 _365_/Q _237_/Q VGND VGND VPWR VPWR final_adder.U$$187/B1 final_adder.U$$186/B
+ sky130_fd_sc_hd__ha_1
XU$$3298 U$$3846/A1 U$$3340/A2 U$$3298/B1 U$$3340/B2 VGND VGND VPWR VPWR U$$3299/A
+ sky130_fd_sc_hd__a22o_1
XU$$2553 U$$2553/A U$$2591/B VGND VGND VPWR VPWR U$$2553/X sky130_fd_sc_hd__xor2_1
XU$$2564 U$$2973/B1 U$$2574/A2 U$$2840/A1 U$$2574/B2 VGND VGND VPWR VPWR U$$2565/A
+ sky130_fd_sc_hd__a22o_1
XU$$1830 U$$1830/A U$$1832/B VGND VGND VPWR VPWR U$$1830/X sky130_fd_sc_hd__xor2_1
XU$$2575 U$$2575/A U$$2575/B VGND VGND VPWR VPWR U$$2575/X sky130_fd_sc_hd__xor2_1
XU$$2586 U$$4365/B1 U$$2598/A2 U$$4367/B1 U$$2598/B2 VGND VGND VPWR VPWR U$$2587/A
+ sky130_fd_sc_hd__a22o_1
XU$$1841 U$$882/A1 U$$1841/A2 U$$882/B1 U$$1841/B2 VGND VGND VPWR VPWR U$$1842/A sky130_fd_sc_hd__a22o_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1852 U$$1852/A U$$1854/B VGND VGND VPWR VPWR U$$1852/X sky130_fd_sc_hd__xor2_1
XU$$2597 U$$2597/A U$$2602/A VGND VGND VPWR VPWR U$$2597/X sky130_fd_sc_hd__xor2_1
XU$$1863 U$$3370/A1 U$$1909/A2 U$$3370/B1 U$$1909/B2 VGND VGND VPWR VPWR U$$1864/A
+ sky130_fd_sc_hd__a22o_1
XU$$1874 U$$1874/A U$$1874/B VGND VGND VPWR VPWR U$$1874/X sky130_fd_sc_hd__xor2_1
XU$$1885 U$$4486/B1 U$$1915/A2 U$$4353/A1 U$$1915/B2 VGND VGND VPWR VPWR U$$1886/A
+ sky130_fd_sc_hd__a22o_1
XU$$1896 U$$1896/A U$$1918/A VGND VGND VPWR VPWR U$$1896/X sky130_fd_sc_hd__xor2_1
XFILLER_148_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_97_0 dadda_fa_5_97_0/A dadda_fa_5_97_0/B dadda_fa_5_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_98_0/A dadda_fa_6_97_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_174_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$515 final_adder.U$$514/B final_adder.U$$399/X final_adder.U$$391/X
+ VGND VGND VPWR VPWR final_adder.U$$515/X sky130_fd_sc_hd__a21o_1
XFILLER_84_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$526 final_adder.U$$534/B final_adder.U$$526/B VGND VGND VPWR VPWR
+ final_adder.U$$646/B sky130_fd_sc_hd__and2_1
XFILLER_57_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$537 final_adder.U$$536/B final_adder.U$$421/X final_adder.U$$413/X
+ VGND VGND VPWR VPWR final_adder.U$$537/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$548 final_adder.U$$556/B final_adder.U$$548/B VGND VGND VPWR VPWR
+ final_adder.U$$668/B sky130_fd_sc_hd__and2_1
XFILLER_85_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$559 final_adder.U$$558/B final_adder.U$$443/X final_adder.U$$435/X
+ VGND VGND VPWR VPWR final_adder.U$$559/X sky130_fd_sc_hd__a21o_1
XFILLER_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$409 U$$409/A U$$410/A VGND VGND VPWR VPWR U$$409/X sky130_fd_sc_hd__xor2_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_106_1 U$$3943/X U$$4076/X U$$4209/X VGND VGND VPWR VPWR dadda_fa_4_107_0/CIN
+ dadda_fa_4_106_2/A sky130_fd_sc_hd__fa_1
XFILLER_106_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_127_0 U$$4383/Y U$$4517/X input159/X VGND VGND VPWR VPWR dadda_fa_6_127_0/COUT
+ dadda_fa_7_127_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_47_3 dadda_fa_3_47_3/A dadda_fa_3_47_3/B dadda_fa_3_47_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_1/B dadda_fa_4_47_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_75_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$910 U$$910/A1 U$$910/A2 U$$912/A1 U$$910/B2 VGND VGND VPWR VPWR U$$911/A sky130_fd_sc_hd__a22o_1
XU$$921 U$$921/A U$$958/A VGND VGND VPWR VPWR U$$921/X sky130_fd_sc_hd__xor2_1
XFILLER_29_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$932 U$$932/A1 U$$942/A2 U$$934/A1 U$$942/B2 VGND VGND VPWR VPWR U$$933/A sky130_fd_sc_hd__a22o_1
XU$$943 U$$943/A U$$943/B VGND VGND VPWR VPWR U$$943/X sky130_fd_sc_hd__xor2_1
XFILLER_28_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$954 U$$954/A1 U$$956/A2 U$$956/A1 U$$956/B2 VGND VGND VPWR VPWR U$$955/A sky130_fd_sc_hd__a22o_1
XFILLER_62_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1104 U$$967/A1 U$$1170/A2 U$$969/A1 U$$1170/B2 VGND VGND VPWR VPWR U$$1105/A sky130_fd_sc_hd__a22o_1
XU$$965 U$$965/A1 U$$979/A2 U$$965/B1 U$$979/B2 VGND VGND VPWR VPWR U$$966/A sky130_fd_sc_hd__a22o_1
XU$$1115 U$$1115/A U$$1171/B VGND VGND VPWR VPWR U$$1115/X sky130_fd_sc_hd__xor2_1
XU$$976 U$$976/A U$$980/B VGND VGND VPWR VPWR U$$976/X sky130_fd_sc_hd__xor2_1
XU$$1126 U$$989/A1 U$$1164/A2 U$$991/A1 U$$1164/B2 VGND VGND VPWR VPWR U$$1127/A sky130_fd_sc_hd__a22o_1
XU$$987 U$$987/A1 U$$999/A2 U$$987/B1 U$$999/B2 VGND VGND VPWR VPWR U$$988/A sky130_fd_sc_hd__a22o_1
XU$$1137 U$$1137/A U$$1175/B VGND VGND VPWR VPWR U$$1137/X sky130_fd_sc_hd__xor2_1
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$998 U$$998/A U$$998/B VGND VGND VPWR VPWR U$$998/X sky130_fd_sc_hd__xor2_1
XU$$1148 U$$50/B1 U$$1170/A2 U$$739/A1 U$$1170/B2 VGND VGND VPWR VPWR U$$1149/A sky130_fd_sc_hd__a22o_1
XU$$1159 U$$1159/A U$$1163/B VGND VGND VPWR VPWR U$$1159/X sky130_fd_sc_hd__xor2_1
XFILLER_102_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1260 input62/X VGND VGND VPWR VPWR U$$547/A sky130_fd_sc_hd__buf_6
Xfanout1271 fanout1279/X VGND VGND VPWR VPWR U$$4159/B sky130_fd_sc_hd__buf_4
Xfanout1282 U$$407/B VGND VGND VPWR VPWR U$$411/A sky130_fd_sc_hd__buf_4
Xfanout1293 fanout1299/X VGND VGND VPWR VPWR U$$4110/A sky130_fd_sc_hd__buf_4
Xdadda_fa_2_42_2 U$$2751/X U$$2884/X U$$2926/B VGND VGND VPWR VPWR dadda_fa_3_43_1/A
+ dadda_fa_3_42_3/A sky130_fd_sc_hd__fa_1
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3040 U$$4410/A1 U$$3122/A2 U$$4412/A1 U$$3122/B2 VGND VGND VPWR VPWR U$$3041/A
+ sky130_fd_sc_hd__a22o_1
XU$$3051 U$$3051/A U$$3073/B VGND VGND VPWR VPWR U$$3051/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_35_1 U$$742/X U$$875/X U$$1008/X VGND VGND VPWR VPWR dadda_fa_3_36_0/CIN
+ dadda_fa_3_35_2/CIN sky130_fd_sc_hd__fa_1
XU$$3062 U$$4158/A1 U$$3072/A2 U$$4295/B1 U$$3072/B2 VGND VGND VPWR VPWR U$$3063/A
+ sky130_fd_sc_hd__a22o_1
XU$$3073 U$$3073/A U$$3073/B VGND VGND VPWR VPWR U$$3073/X sky130_fd_sc_hd__xor2_1
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3084 U$$4454/A1 U$$3148/A2 U$$4456/A1 U$$3148/B2 VGND VGND VPWR VPWR U$$3085/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_12_0 input160/X dadda_fa_5_12_0/B dadda_fa_5_12_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_6_13_0/A dadda_fa_6_12_0/CIN sky130_fd_sc_hd__fa_1
XU$$3095 U$$3095/A U$$3107/B VGND VGND VPWR VPWR U$$3095/X sky130_fd_sc_hd__xor2_1
XU$$2350 U$$2350/A U$$2402/B VGND VGND VPWR VPWR U$$2350/X sky130_fd_sc_hd__xor2_1
XU$$2361 U$$989/B1 U$$2395/A2 U$$856/A1 U$$2395/B2 VGND VGND VPWR VPWR U$$2362/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_28_0 U$$63/X U$$196/X U$$329/X VGND VGND VPWR VPWR dadda_fa_3_29_1/CIN
+ dadda_fa_3_28_3/A sky130_fd_sc_hd__fa_1
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2372 U$$2372/A U$$2416/B VGND VGND VPWR VPWR U$$2372/X sky130_fd_sc_hd__xor2_1
XU$$2383 U$$876/A1 U$$2415/A2 U$$878/A1 U$$2415/B2 VGND VGND VPWR VPWR U$$2384/A sky130_fd_sc_hd__a22o_1
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2394 U$$2394/A U$$2396/B VGND VGND VPWR VPWR U$$2394/X sky130_fd_sc_hd__xor2_1
XU$$1660 U$$2891/B1 U$$1696/A2 U$$2758/A1 U$$1696/B2 VGND VGND VPWR VPWR U$$1661/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1671 U$$1671/A U$$1703/B VGND VGND VPWR VPWR U$$1671/X sky130_fd_sc_hd__xor2_1
XFILLER_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1682 U$$721/B1 U$$1698/A2 U$$999/A1 U$$1698/B2 VGND VGND VPWR VPWR U$$1683/A sky130_fd_sc_hd__a22o_1
XU$$1693 U$$1693/A U$$1697/B VGND VGND VPWR VPWR U$$1693/X sky130_fd_sc_hd__xor2_1
XFILLER_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_87_4 U$$3240/X U$$3373/X U$$3506/X VGND VGND VPWR VPWR dadda_fa_2_88_4/B
+ dadda_fa_3_87_0/A sky130_fd_sc_hd__fa_1
XFILLER_118_1013 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_57_2 dadda_fa_4_57_2/A dadda_fa_4_57_2/B dadda_fa_4_57_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_58_0/CIN dadda_fa_5_57_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$301 final_adder.U$$300/B final_adder.U$$175/X final_adder.U$$173/X
+ VGND VGND VPWR VPWR final_adder.U$$301/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$312 final_adder.U$$314/B final_adder.U$$312/B VGND VGND VPWR VPWR
+ final_adder.U$$438/B sky130_fd_sc_hd__and2_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$323 final_adder.U$$322/B final_adder.U$$197/X final_adder.U$$195/X
+ VGND VGND VPWR VPWR final_adder.U$$323/X sky130_fd_sc_hd__a21o_1
XFILLER_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$334 final_adder.U$$336/B final_adder.U$$334/B VGND VGND VPWR VPWR
+ final_adder.U$$460/B sky130_fd_sc_hd__and2_1
XFILLER_58_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$345 final_adder.U$$344/B final_adder.U$$219/X final_adder.U$$217/X
+ VGND VGND VPWR VPWR final_adder.U$$345/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$356 final_adder.U$$358/B final_adder.U$$356/B VGND VGND VPWR VPWR
+ final_adder.U$$482/B sky130_fd_sc_hd__and2_1
Xdadda_fa_7_27_0 dadda_fa_7_27_0/A dadda_fa_7_27_0/B dadda_fa_7_27_0/CIN VGND VGND
+ VPWR VPWR _324_/D _195_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$367 final_adder.U$$366/B final_adder.U$$241/X final_adder.U$$239/X
+ VGND VGND VPWR VPWR final_adder.U$$367/X sky130_fd_sc_hd__a21o_1
XU$$206 U$$206/A U$$210/B VGND VGND VPWR VPWR U$$206/X sky130_fd_sc_hd__xor2_1
XFILLER_85_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$378 final_adder.U$$378/A final_adder.U$$378/B VGND VGND VPWR VPWR
+ final_adder.U$$500/A sky130_fd_sc_hd__and2_1
XU$$217 U$$902/A1 U$$219/A2 U$$902/B1 U$$219/B2 VGND VGND VPWR VPWR U$$218/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$389 final_adder.U$$388/B final_adder.U$$267/X final_adder.U$$263/X
+ VGND VGND VPWR VPWR final_adder.U$$389/X sky130_fd_sc_hd__a21o_1
XU$$228 U$$228/A U$$230/B VGND VGND VPWR VPWR U$$228/X sky130_fd_sc_hd__xor2_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$239 U$$787/A1 U$$253/A2 U$$787/B1 U$$253/B2 VGND VGND VPWR VPWR U$$240/A sky130_fd_sc_hd__a22o_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_52_1 dadda_fa_3_52_1/A dadda_fa_3_52_1/B dadda_fa_3_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_0/CIN dadda_fa_4_52_2/A sky130_fd_sc_hd__fa_1
XFILLER_48_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_68_1 U$$675/X U$$808/X U$$941/X VGND VGND VPWR VPWR dadda_fa_1_69_6/A
+ dadda_fa_1_68_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_45_0 dadda_fa_3_45_0/A dadda_fa_3_45_0/B dadda_fa_3_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_0/B dadda_fa_4_45_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$740 U$$740/A U$$744/B VGND VGND VPWR VPWR U$$740/X sky130_fd_sc_hd__xor2_1
XU$$751 U$$66/A1 U$$769/A2 U$$68/A1 U$$769/B2 VGND VGND VPWR VPWR U$$752/A sky130_fd_sc_hd__a22o_1
XU$$762 U$$762/A U$$764/B VGND VGND VPWR VPWR U$$762/X sky130_fd_sc_hd__xor2_1
XU$$773 U$$773/A1 U$$817/A2 U$$773/B1 U$$817/B2 VGND VGND VPWR VPWR U$$774/A sky130_fd_sc_hd__a22o_1
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$784 U$$784/A U$$820/B VGND VGND VPWR VPWR U$$784/X sky130_fd_sc_hd__xor2_1
XU$$795 U$$932/A1 U$$809/A2 U$$934/A1 U$$809/B2 VGND VGND VPWR VPWR U$$796/A sky130_fd_sc_hd__a22o_1
XFILLER_31_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_2_98_5 U$$4326/X U$$4459/X VGND VGND VPWR VPWR dadda_fa_3_99_2/B dadda_fa_4_98_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_31_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_102_0 dadda_fa_7_102_0/A dadda_fa_7_102_0/B dadda_fa_7_102_0/CIN VGND
+ VGND VPWR VPWR _399_/D _270_/D sky130_fd_sc_hd__fa_1
XFILLER_144_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_97_3 U$$3526/X U$$3659/X U$$3792/X VGND VGND VPWR VPWR dadda_fa_3_98_1/B
+ dadda_fa_3_97_3/B sky130_fd_sc_hd__fa_1
XFILLER_160_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_67_1 dadda_fa_5_67_1/A dadda_fa_5_67_1/B dadda_fa_5_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_68_0/B dadda_fa_7_67_0/A sky130_fd_sc_hd__fa_1
XFILLER_4_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_867 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout508 U$$3251/A2 VGND VGND VPWR VPWR U$$3285/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout519 U$$3018/X VGND VGND VPWR VPWR U$$3118/A2 sky130_fd_sc_hd__buf_4
XFILLER_101_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_59_8 dadda_fa_1_59_8/A dadda_fa_1_59_8/B dadda_fa_1_59_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_60_3/A dadda_fa_3_59_0/A sky130_fd_sc_hd__fa_2
XFILLER_82_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1090 input82/X VGND VGND VPWR VPWR U$$878/B1 sky130_fd_sc_hd__buf_6
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_106_0 dadda_fa_2_106_0/A U$$3012/X U$$3145/X VGND VGND VPWR VPWR dadda_fa_3_107_3/B
+ dadda_fa_3_106_3/CIN sky130_fd_sc_hd__fa_1
XU$$2180 U$$2180/A U$$2186/B VGND VGND VPWR VPWR U$$2180/X sky130_fd_sc_hd__xor2_1
XU$$2191 U$$2191/A VGND VGND VPWR VPWR U$$2191/Y sky130_fd_sc_hd__inv_1
XFILLER_50_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1490 U$$120/A1 U$$1502/A2 U$$120/B1 U$$1502/B2 VGND VGND VPWR VPWR U$$1491/A sky130_fd_sc_hd__a22o_1
XFILLER_22_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_85_1 U$$1906/X U$$2039/X U$$2172/X VGND VGND VPWR VPWR dadda_fa_2_86_2/CIN
+ dadda_fa_2_85_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_62_0 dadda_fa_4_62_0/A dadda_fa_4_62_0/B dadda_fa_4_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_63_0/A dadda_fa_5_62_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_78_0 U$$1227/X U$$1360/X U$$1493/X VGND VGND VPWR VPWR dadda_fa_2_79_0/B
+ dadda_fa_2_78_3/B sky130_fd_sc_hd__fa_1
XFILLER_77_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$120 _416_/Q _288_/Q VGND VGND VPWR VPWR final_adder.U$$905/B1 final_adder.U$$134/A
+ sky130_fd_sc_hd__ha_1
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$131 final_adder.U$$130/B final_adder.U$$901/B1 final_adder.U$$131/B1
+ VGND VGND VPWR VPWR final_adder.U$$131/X sky130_fd_sc_hd__a21o_1
XU$$3809 U$$4492/B1 U$$3833/A2 U$$4359/A1 U$$3833/B2 VGND VGND VPWR VPWR U$$3810/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$142 final_adder.U$$142/A final_adder.U$$142/B VGND VGND VPWR VPWR
+ final_adder.U$$270/B sky130_fd_sc_hd__and2_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$153 final_adder.U$$152/B final_adder.U$$923/B1 final_adder.U$$153/B1
+ VGND VGND VPWR VPWR final_adder.U$$153/X sky130_fd_sc_hd__a21o_1
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$164 final_adder.U$$164/A final_adder.U$$164/B VGND VGND VPWR VPWR
+ final_adder.U$$292/B sky130_fd_sc_hd__and2_1
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$175 final_adder.U$$174/B final_adder.U$$945/B1 final_adder.U$$175/B1
+ VGND VGND VPWR VPWR final_adder.U$$175/X sky130_fd_sc_hd__a21o_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$186 final_adder.U$$186/A final_adder.U$$186/B VGND VGND VPWR VPWR
+ final_adder.U$$314/B sky130_fd_sc_hd__and2_1
XFILLER_73_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$197 final_adder.U$$196/B final_adder.U$$967/B1 final_adder.U$$197/B1
+ VGND VGND VPWR VPWR final_adder.U$$197/X sky130_fd_sc_hd__a21o_1
XFILLER_73_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_383_ _383_/CLK _383_/D VGND VGND VPWR VPWR _383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_77_0 dadda_fa_6_77_0/A dadda_fa_6_77_0/B dadda_fa_6_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_78_0/B dadda_fa_7_77_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput160 c[12] VGND VGND VPWR VPWR input160/X sky130_fd_sc_hd__clkbuf_4
Xinput171 c[22] VGND VGND VPWR VPWR input171/X sky130_fd_sc_hd__buf_2
Xinput182 c[32] VGND VGND VPWR VPWR input182/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput193 c[42] VGND VGND VPWR VPWR input193/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$570 U$$707/A1 U$$638/A2 U$$709/A1 U$$638/B2 VGND VGND VPWR VPWR U$$571/A sky130_fd_sc_hd__a22o_1
XFILLER_17_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$581 U$$581/A U$$607/B VGND VGND VPWR VPWR U$$581/X sky130_fd_sc_hd__xor2_1
XU$$592 U$$864/B1 U$$630/A2 U$$729/B1 U$$630/B2 VGND VGND VPWR VPWR U$$593/A sky130_fd_sc_hd__a22o_1
XFILLER_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_95_0 U$$2591/X U$$2724/X U$$2857/X VGND VGND VPWR VPWR dadda_fa_3_96_0/B
+ dadda_fa_3_95_2/B sky130_fd_sc_hd__fa_1
XFILLER_173_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_71_7 dadda_fa_1_71_7/A dadda_fa_1_71_7/B dadda_fa_1_71_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_72_2/CIN dadda_fa_2_71_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_115_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_6 dadda_fa_1_64_6/A dadda_fa_1_64_6/B dadda_fa_1_64_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_65_2/B dadda_fa_2_64_5/B sky130_fd_sc_hd__fa_1
XFILLER_101_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_57_5 U$$3180/X U$$3313/X U$$3446/X VGND VGND VPWR VPWR dadda_fa_2_58_2/A
+ dadda_fa_2_57_5/A sky130_fd_sc_hd__fa_1
XFILLER_28_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1028 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_94_0 dadda_fa_7_94_0/A dadda_fa_7_94_0/B dadda_fa_7_94_0/CIN VGND VGND
+ VPWR VPWR _391_/D _262_/D sky130_fd_sc_hd__fa_1
XFILLER_149_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout850 U$$2052/B2 VGND VGND VPWR VPWR U$$2044/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout861 U$$1786/X VGND VGND VPWR VPWR U$$1891/B2 sky130_fd_sc_hd__buf_6
XU$$4307 U$$4307/A1 U$$4381/A2 U$$4307/B1 U$$4381/B2 VGND VGND VPWR VPWR U$$4308/A
+ sky130_fd_sc_hd__a22o_1
Xfanout872 U$$1593/B2 VGND VGND VPWR VPWR U$$1567/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4318 U$$4318/A U$$4350/B VGND VGND VPWR VPWR U$$4318/X sky130_fd_sc_hd__xor2_1
Xfanout883 U$$142/X VGND VGND VPWR VPWR U$$259/B2 sky130_fd_sc_hd__clkbuf_8
XU$$4329 U$$4464/B1 U$$4349/A2 U$$4331/A1 U$$4349/B2 VGND VGND VPWR VPWR U$$4330/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout894 U$$1480/B2 VGND VGND VPWR VPWR U$$1502/B2 sky130_fd_sc_hd__buf_6
XU$$3606 U$$4152/B1 U$$3644/A2 U$$4017/B1 U$$3644/B2 VGND VGND VPWR VPWR U$$3607/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3617 U$$3617/A U$$3695/B VGND VGND VPWR VPWR U$$3617/X sky130_fd_sc_hd__xor2_1
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3628 U$$3628/A1 U$$3640/A2 U$$3628/B1 U$$3640/B2 VGND VGND VPWR VPWR U$$3629/A
+ sky130_fd_sc_hd__a22o_1
XU$$3639 U$$3639/A U$$3641/B VGND VGND VPWR VPWR U$$3639/X sky130_fd_sc_hd__xor2_1
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2905 U$$3314/B1 U$$2989/A2 U$$3181/A1 U$$2989/B2 VGND VGND VPWR VPWR U$$2906/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2916 U$$2916/A U$$2944/B VGND VGND VPWR VPWR U$$2916/X sky130_fd_sc_hd__xor2_1
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2927 U$$3338/A1 U$$2937/A2 U$$735/B1 U$$2937/B2 VGND VGND VPWR VPWR U$$2928/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2938 U$$2938/A U$$2938/B VGND VGND VPWR VPWR U$$2938/X sky130_fd_sc_hd__xor2_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_22_2 U$$1115/X U$$1248/X U$$1381/X VGND VGND VPWR VPWR dadda_fa_4_23_1/A
+ dadda_fa_4_22_2/B sky130_fd_sc_hd__fa_1
XU$$2949 U$$4456/A1 U$$3005/A2 U$$4456/B1 U$$3005/B2 VGND VGND VPWR VPWR U$$2950/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_366_ _366_/CLK _366_/D VGND VGND VPWR VPWR _366_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_174_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_297_ _319_/CLK _297_/D VGND VGND VPWR VPWR _297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_74_5 dadda_fa_2_74_5/A dadda_fa_2_74_5/B dadda_fa_2_74_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_2/A dadda_fa_4_74_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_67_4 dadda_fa_2_67_4/A dadda_fa_2_67_4/B dadda_fa_2_67_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_1/CIN dadda_fa_3_67_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$0_1780 VGND VGND VPWR VPWR U$$0_1780/HI U$$0/A sky130_fd_sc_hd__conb_1
XFILLER_24_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4421_1858 VGND VGND VPWR VPWR U$$4421_1858/HI U$$4421/B sky130_fd_sc_hd__conb_1
XFILLER_137_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_104_1 dadda_fa_5_104_1/A dadda_fa_5_104_1/B dadda_fa_5_104_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_105_0/B dadda_fa_7_104_0/A sky130_fd_sc_hd__fa_1
XFILLER_172_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_62_3 U$$3589/X U$$3722/X U$$3855/X VGND VGND VPWR VPWR dadda_fa_2_63_1/B
+ dadda_fa_2_62_4/B sky130_fd_sc_hd__fa_1
XFILLER_47_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_55_2 U$$1580/X U$$1713/X U$$1846/X VGND VGND VPWR VPWR dadda_fa_2_56_1/A
+ dadda_fa_2_55_4/A sky130_fd_sc_hd__fa_1
XFILLER_67_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1367_1786 VGND VGND VPWR VPWR U$$1367_1786/HI U$$1367/B1 sky130_fd_sc_hd__conb_1
Xdadda_fa_4_32_1 dadda_fa_4_32_1/A dadda_fa_4_32_1/B dadda_fa_4_32_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_33_0/B dadda_fa_5_32_1/B sky130_fd_sc_hd__fa_1
XFILLER_83_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_48_1 U$$502/X U$$635/X U$$768/X VGND VGND VPWR VPWR dadda_fa_2_49_1/B
+ dadda_fa_2_48_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_25_0 dadda_fa_4_25_0/A dadda_fa_4_25_0/B dadda_fa_4_25_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_26_0/A dadda_fa_5_25_1/A sky130_fd_sc_hd__fa_1
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_220_ _349_/CLK _220_/D VGND VGND VPWR VPWR _220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_77_3 dadda_fa_3_77_3/A dadda_fa_3_77_3/B dadda_fa_3_77_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_1/B dadda_fa_4_77_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_151_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1601 U$$2042/A1 VGND VGND VPWR VPWR U$$672/A1 sky130_fd_sc_hd__buf_4
XFILLER_104_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1612 U$$2860/B1 VGND VGND VPWR VPWR U$$2175/B1 sky130_fd_sc_hd__buf_6
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1623 U$$4504/A1 VGND VGND VPWR VPWR U$$4365/B1 sky130_fd_sc_hd__buf_4
Xfanout1634 U$$4502/A1 VGND VGND VPWR VPWR U$$4226/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1645 input114/X VGND VGND VPWR VPWR U$$4500/A1 sky130_fd_sc_hd__buf_2
Xfanout1656 U$$2578/A1 VGND VGND VPWR VPWR U$$2576/B1 sky130_fd_sc_hd__buf_6
XU$$4104 U$$4104/A U$$4108/B VGND VGND VPWR VPWR U$$4104/X sky130_fd_sc_hd__xor2_1
XU$$4115 U$$4113/B U$$4110/A input57/X U$$4110/Y VGND VGND VPWR VPWR U$$4115/X sky130_fd_sc_hd__a22o_2
Xfanout1667 U$$4494/A1 VGND VGND VPWR VPWR U$$384/A1 sky130_fd_sc_hd__buf_2
Xfanout680 U$$638/B2 VGND VGND VPWR VPWR U$$610/B2 sky130_fd_sc_hd__buf_4
XU$$4126 U$$4400/A1 U$$4158/A2 U$$4400/B1 U$$4158/B2 VGND VGND VPWR VPWR U$$4127/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1678 fanout1680/X VGND VGND VPWR VPWR U$$4492/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1689 U$$1358/B VGND VGND VPWR VPWR U$$1364/B sky130_fd_sc_hd__buf_6
XU$$4137 U$$4137/A U$$4159/B VGND VGND VPWR VPWR U$$4137/X sky130_fd_sc_hd__xor2_1
Xfanout691 U$$4309/B2 VGND VGND VPWR VPWR U$$4325/B2 sky130_fd_sc_hd__buf_6
XU$$3403 U$$3403/A U$$3411/B VGND VGND VPWR VPWR U$$3403/X sky130_fd_sc_hd__xor2_1
XFILLER_93_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_3_14_0 U$$35/X U$$168/X VGND VGND VPWR VPWR dadda_fa_4_15_2/B dadda_ha_3_14_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$4148 U$$4422/A1 U$$4240/A2 U$$4150/A1 U$$4240/B2 VGND VGND VPWR VPWR U$$4149/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4159 U$$4159/A U$$4159/B VGND VGND VPWR VPWR U$$4159/X sky130_fd_sc_hd__xor2_1
XU$$3414 U$$3551/A1 U$$3416/A2 U$$3416/A1 U$$3416/B2 VGND VGND VPWR VPWR U$$3415/A
+ sky130_fd_sc_hd__a22o_1
XU$$3425 U$$3425/A VGND VGND VPWR VPWR U$$3425/Y sky130_fd_sc_hd__inv_1
XFILLER_18_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3436 U$$3436/A U$$3482/B VGND VGND VPWR VPWR U$$3436/X sky130_fd_sc_hd__xor2_1
XU$$2702 U$$2702/A U$$2708/B VGND VGND VPWR VPWR U$$2702/X sky130_fd_sc_hd__xor2_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3447 U$$707/A1 U$$3523/A2 U$$3447/B1 U$$3523/B2 VGND VGND VPWR VPWR U$$3448/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3458 U$$3458/A U$$3468/B VGND VGND VPWR VPWR U$$3458/X sky130_fd_sc_hd__xor2_1
XU$$2713 U$$4220/A1 U$$2733/A2 U$$4220/B1 U$$2733/B2 VGND VGND VPWR VPWR U$$2714/A
+ sky130_fd_sc_hd__a22o_1
XU$$2724 U$$2724/A U$$2724/B VGND VGND VPWR VPWR U$$2724/X sky130_fd_sc_hd__xor2_1
XU$$3469 U$$4428/A1 U$$3471/A2 U$$4291/B1 U$$3471/B2 VGND VGND VPWR VPWR U$$3470/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2735 U$$3418/B1 U$$2737/A2 U$$3285/A1 U$$2737/B2 VGND VGND VPWR VPWR U$$2736/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2746 U$$2746/A1 U$$2804/A2 U$$2748/A1 U$$2804/B2 VGND VGND VPWR VPWR U$$2747/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2757 U$$2757/A U$$2799/B VGND VGND VPWR VPWR U$$2757/X sky130_fd_sc_hd__xor2_1
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2768 U$$3314/B1 U$$2856/A2 U$$30/A1 U$$2856/B2 VGND VGND VPWR VPWR U$$2769/A sky130_fd_sc_hd__a22o_1
XFILLER_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2779 U$$2779/A U$$2811/B VGND VGND VPWR VPWR U$$2779/X sky130_fd_sc_hd__xor2_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_418_ _421_/CLK _418_/D VGND VGND VPWR VPWR _418_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_349_ _349_/CLK _349_/D VGND VGND VPWR VPWR _349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_72_2 dadda_fa_2_72_2/A dadda_fa_2_72_2/B dadda_fa_2_72_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_1/A dadda_fa_3_72_3/A sky130_fd_sc_hd__fa_1
XFILLER_130_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_65_1 dadda_fa_2_65_1/A dadda_fa_2_65_1/B dadda_fa_2_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_0/CIN dadda_fa_3_65_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_97_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$708 final_adder.U$$708/A final_adder.U$$708/B VGND VGND VPWR VPWR
+ final_adder.U$$788/A sky130_fd_sc_hd__and2_1
XFILLER_110_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$719 final_adder.U$$718/B final_adder.U$$615/X final_adder.U$$599/X
+ VGND VGND VPWR VPWR final_adder.U$$719/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_5_42_0 dadda_fa_5_42_0/A dadda_fa_5_42_0/B dadda_fa_5_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_43_0/A dadda_fa_6_42_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_58_0 dadda_fa_2_58_0/A dadda_fa_2_58_0/B dadda_fa_2_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_0/B dadda_fa_3_58_2/B sky130_fd_sc_hd__fa_1
XFILLER_56_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3970 U$$4107/A1 U$$3970/A2 U$$3970/B1 U$$3970/B2 VGND VGND VPWR VPWR U$$3971/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3981 U$$3981/A1 U$$4005/A2 U$$4257/A1 U$$4005/B2 VGND VGND VPWR VPWR U$$3982/A
+ sky130_fd_sc_hd__a22o_1
XU$$3992 U$$3992/A U$$4026/B VGND VGND VPWR VPWR U$$3992/X sky130_fd_sc_hd__xor2_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_87_2 dadda_fa_4_87_2/A dadda_fa_4_87_2/B dadda_fa_4_87_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_88_0/CIN dadda_fa_5_87_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_146_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput261 output261/A VGND VGND VPWR VPWR o[103] sky130_fd_sc_hd__buf_2
Xdadda_fa_7_57_0 dadda_fa_7_57_0/A dadda_fa_7_57_0/B dadda_fa_7_57_0/CIN VGND VGND
+ VPWR VPWR _354_/D _225_/D sky130_fd_sc_hd__fa_1
Xoutput272 output272/A VGND VGND VPWR VPWR o[113] sky130_fd_sc_hd__buf_2
Xoutput283 output283/A VGND VGND VPWR VPWR o[123] sky130_fd_sc_hd__buf_2
Xoutput294 output294/A VGND VGND VPWR VPWR o[18] sky130_fd_sc_hd__buf_2
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_60_0 U$$1989/X U$$2122/X U$$2255/X VGND VGND VPWR VPWR dadda_fa_2_61_0/B
+ dadda_fa_2_60_3/B sky130_fd_sc_hd__fa_1
XFILLER_87_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1230_1783 VGND VGND VPWR VPWR U$$1230_1783/HI U$$1230/B1 sky130_fd_sc_hd__conb_1
XFILLER_75_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2009 U$$2009/A U$$2053/B VGND VGND VPWR VPWR U$$2009/X sky130_fd_sc_hd__xor2_1
XFILLER_55_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1308 U$$1308/A U$$1320/B VGND VGND VPWR VPWR U$$1308/X sky130_fd_sc_hd__xor2_1
XU$$1319 U$$906/B1 U$$1359/A2 U$$773/A1 U$$1359/B2 VGND VGND VPWR VPWR U$$1320/A sky130_fd_sc_hd__a22o_1
XFILLER_15_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_203_ _344_/CLK _203_/D VGND VGND VPWR VPWR _203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1102 final_adder.U$$176/A final_adder.U$$885/X VGND VGND VPWR VPWR
+ output360/A sky130_fd_sc_hd__xor2_1
XFILLER_7_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1113 final_adder.U$$166/B final_adder.U$$937/X VGND VGND VPWR VPWR
+ output372/A sky130_fd_sc_hd__xor2_1
XFILLER_23_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1124 final_adder.U$$154/A final_adder.U$$863/X VGND VGND VPWR VPWR
+ output258/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1135 final_adder.U$$144/B final_adder.U$$915/X VGND VGND VPWR VPWR
+ output270/A sky130_fd_sc_hd__xor2_1
XFILLER_7_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1146 final_adder.U$$132/A final_adder.U$$841/X VGND VGND VPWR VPWR
+ output282/A sky130_fd_sc_hd__xor2_1
XFILLER_139_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_82_1 dadda_fa_3_82_1/A dadda_fa_3_82_1/B dadda_fa_3_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_0/CIN dadda_fa_4_82_2/A sky130_fd_sc_hd__fa_1
XFILLER_125_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_75_0 dadda_fa_3_75_0/A dadda_fa_3_75_0/B dadda_fa_3_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_0/B dadda_fa_4_75_1/CIN sky130_fd_sc_hd__fa_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1420 U$$768/B VGND VGND VPWR VPWR U$$764/B sky130_fd_sc_hd__buf_6
XFILLER_79_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1431 U$$2408/B VGND VGND VPWR VPWR U$$2466/A sky130_fd_sc_hd__buf_4
XFILLER_39_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1442 U$$2283/B VGND VGND VPWR VPWR U$$2249/B sky130_fd_sc_hd__clkbuf_4
XFILLER_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1453 input25/X VGND VGND VPWR VPWR U$$2140/B sky130_fd_sc_hd__buf_4
XFILLER_120_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1464 U$$2031/B VGND VGND VPWR VPWR U$$2055/A sky130_fd_sc_hd__buf_2
Xfanout1475 input20/X VGND VGND VPWR VPWR U$$1874/B sky130_fd_sc_hd__buf_6
Xfanout1486 U$$1594/B VGND VGND VPWR VPWR U$$1564/B sky130_fd_sc_hd__buf_6
XU$$3200 U$$3200/A U$$3208/B VGND VGND VPWR VPWR U$$3200/X sky130_fd_sc_hd__xor2_1
Xfanout1497 U$$1461/B VGND VGND VPWR VPWR U$$1433/B sky130_fd_sc_hd__clkbuf_4
XFILLER_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3211 input83/X U$$3255/A2 input84/X U$$3255/B2 VGND VGND VPWR VPWR U$$3212/A sky130_fd_sc_hd__a22o_1
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3222 U$$3222/A U$$3288/A VGND VGND VPWR VPWR U$$3222/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_111_1 dadda_fa_4_111_1/A dadda_fa_4_111_1/B dadda_fa_4_111_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_112_0/B dadda_fa_5_111_1/B sky130_fd_sc_hd__fa_1
XU$$3233 U$$3370/A1 U$$3241/A2 U$$3370/B1 U$$3241/B2 VGND VGND VPWR VPWR U$$3234/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$15 _311_/Q _183_/Q VGND VGND VPWR VPWR final_adder.U$$241/B1 final_adder.U$$240/B
+ sky130_fd_sc_hd__ha_1
XU$$3244 U$$3244/A U$$3288/A VGND VGND VPWR VPWR U$$3244/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$26 _322_/Q _194_/Q VGND VGND VPWR VPWR final_adder.U$$999/B1 final_adder.U$$228/A
+ sky130_fd_sc_hd__ha_1
XU$$2510 U$$4152/B1 U$$2548/A2 U$$4017/B1 U$$2548/B2 VGND VGND VPWR VPWR U$$2511/A
+ sky130_fd_sc_hd__a22o_1
XU$$3255 U$$787/B1 U$$3255/A2 U$$517/A1 U$$3255/B2 VGND VGND VPWR VPWR U$$3256/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$37 _333_/Q _205_/Q VGND VGND VPWR VPWR final_adder.U$$219/B1 final_adder.U$$218/B
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_4_104_0 dadda_fa_4_104_0/A dadda_fa_4_104_0/B dadda_fa_4_104_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_105_0/A dadda_fa_5_104_1/A sky130_fd_sc_hd__fa_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_37_5 dadda_fa_2_37_5/A dadda_fa_2_37_5/B dadda_fa_2_37_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_38_2/A dadda_fa_4_37_0/A sky130_fd_sc_hd__fa_1
XU$$3266 U$$3266/A U$$3284/B VGND VGND VPWR VPWR U$$3266/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$48 _344_/Q _216_/Q VGND VGND VPWR VPWR final_adder.U$$977/B1 final_adder.U$$206/A
+ sky130_fd_sc_hd__ha_1
XFILLER_19_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2521 U$$2521/A U$$2541/B VGND VGND VPWR VPWR U$$2521/X sky130_fd_sc_hd__xor2_1
XU$$2532 U$$66/A1 U$$2532/A2 U$$68/A1 U$$2532/B2 VGND VGND VPWR VPWR U$$2533/A sky130_fd_sc_hd__a22o_1
XFILLER_62_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3277 U$$3551/A1 U$$3285/A2 U$$3416/A1 U$$3285/B2 VGND VGND VPWR VPWR U$$3278/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$59 _355_/Q _227_/Q VGND VGND VPWR VPWR final_adder.U$$197/B1 final_adder.U$$196/B
+ sky130_fd_sc_hd__ha_1
XU$$3288 U$$3288/A VGND VGND VPWR VPWR U$$3288/Y sky130_fd_sc_hd__inv_1
XU$$2543 U$$2543/A U$$2591/B VGND VGND VPWR VPWR U$$2543/X sky130_fd_sc_hd__xor2_1
XU$$3299 U$$3299/A U$$3341/B VGND VGND VPWR VPWR U$$3299/X sky130_fd_sc_hd__xor2_1
XU$$2554 U$$4196/B1 U$$2598/A2 U$$4198/B1 U$$2598/B2 VGND VGND VPWR VPWR U$$2555/A
+ sky130_fd_sc_hd__a22o_1
XU$$1820 U$$1820/A U$$1828/B VGND VGND VPWR VPWR U$$1820/X sky130_fd_sc_hd__xor2_1
XU$$2565 U$$2565/A U$$2575/B VGND VGND VPWR VPWR U$$2565/X sky130_fd_sc_hd__xor2_1
XFILLER_55_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1831 U$$735/A1 U$$1831/A2 U$$52/A1 U$$1831/B2 VGND VGND VPWR VPWR U$$1832/A sky130_fd_sc_hd__a22o_1
XFILLER_22_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2576 U$$2576/A1 U$$2578/A2 U$$2576/B1 U$$2578/B2 VGND VGND VPWR VPWR U$$2577/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2587 U$$2587/A U$$2591/B VGND VGND VPWR VPWR U$$2587/X sky130_fd_sc_hd__xor2_1
XU$$1842 U$$1842/A U$$1854/B VGND VGND VPWR VPWR U$$1842/X sky130_fd_sc_hd__xor2_1
XU$$2598 U$$3418/B1 U$$2598/A2 U$$3285/A1 U$$2598/B2 VGND VGND VPWR VPWR U$$2599/A
+ sky130_fd_sc_hd__a22o_1
XU$$1853 U$$346/A1 U$$1891/A2 U$$2814/A1 U$$1891/B2 VGND VGND VPWR VPWR U$$1854/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1864 U$$1864/A U$$1874/B VGND VGND VPWR VPWR U$$1864/X sky130_fd_sc_hd__xor2_1
XU$$1875 U$$3382/A1 U$$1915/A2 U$$3382/B1 U$$1915/B2 VGND VGND VPWR VPWR U$$1876/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1886 U$$1886/A U$$1916/B VGND VGND VPWR VPWR U$$1886/X sky130_fd_sc_hd__xor2_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1897 U$$2443/B1 U$$1909/A2 U$$2310/A1 U$$1909/B2 VGND VGND VPWR VPWR U$$1898/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_97_1 dadda_fa_5_97_1/A dadda_fa_5_97_1/B dadda_fa_5_97_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_98_0/B dadda_fa_7_97_0/A sky130_fd_sc_hd__fa_1
XFILLER_128_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_980 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$505 final_adder.U$$500/A final_adder.U$$255/X final_adder.U$$379/X
+ VGND VGND VPWR VPWR final_adder.U$$505/X sky130_fd_sc_hd__a21o_2
Xfinal_adder.U$$516 final_adder.U$$524/B final_adder.U$$516/B VGND VGND VPWR VPWR
+ final_adder.U$$636/B sky130_fd_sc_hd__and2_1
XFILLER_29_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$527 final_adder.U$$526/B final_adder.U$$411/X final_adder.U$$403/X
+ VGND VGND VPWR VPWR final_adder.U$$527/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$538 final_adder.U$$546/B final_adder.U$$538/B VGND VGND VPWR VPWR
+ final_adder.U$$658/B sky130_fd_sc_hd__and2_1
XFILLER_57_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$549 final_adder.U$$548/B final_adder.U$$433/X final_adder.U$$425/X
+ VGND VGND VPWR VPWR final_adder.U$$549/X sky130_fd_sc_hd__a21o_1
XFILLER_85_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4490 U$$4490/A1 U$$4388/X U$$4492/A1 U$$4492/B2 VGND VGND VPWR VPWR U$$4491/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_926 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_92_0 dadda_fa_4_92_0/A dadda_fa_4_92_0/B dadda_fa_4_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_93_0/A dadda_fa_5_92_1/A sky130_fd_sc_hd__fa_1
XFILLER_158_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_106_2 U$$4342/X U$$4475/X input136/X VGND VGND VPWR VPWR dadda_fa_4_107_1/A
+ dadda_fa_4_106_2/B sky130_fd_sc_hd__fa_1
XFILLER_134_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4473_1884 VGND VGND VPWR VPWR U$$4473_1884/HI U$$4473/B sky130_fd_sc_hd__conb_1
XFILLER_162_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$900 U$$900/A1 U$$902/A2 U$$900/B1 U$$902/B2 VGND VGND VPWR VPWR U$$901/A sky130_fd_sc_hd__a22o_1
XFILLER_63_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$911 U$$911/A U$$913/B VGND VGND VPWR VPWR U$$911/X sky130_fd_sc_hd__xor2_1
XU$$922 U$$922/A1 U$$952/A2 U$$922/B1 U$$952/B2 VGND VGND VPWR VPWR U$$923/A sky130_fd_sc_hd__a22o_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$933 U$$933/A U$$959/A VGND VGND VPWR VPWR U$$933/X sky130_fd_sc_hd__xor2_1
XFILLER_56_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$944 U$$944/A1 U$$956/A2 U$$944/B1 U$$956/B2 VGND VGND VPWR VPWR U$$945/A sky130_fd_sc_hd__a22o_1
XU$$955 U$$955/A U$$955/B VGND VGND VPWR VPWR U$$955/X sky130_fd_sc_hd__xor2_1
XU$$1105 U$$1105/A U$$1171/B VGND VGND VPWR VPWR U$$1105/X sky130_fd_sc_hd__xor2_1
XFILLER_43_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$966 U$$966/A U$$980/B VGND VGND VPWR VPWR U$$966/X sky130_fd_sc_hd__xor2_1
XU$$1116 U$$2897/A1 U$$1170/A2 U$$2897/B1 U$$1170/B2 VGND VGND VPWR VPWR U$$1117/A
+ sky130_fd_sc_hd__a22o_1
XU$$977 U$$18/A1 U$$979/A2 U$$20/A1 U$$979/B2 VGND VGND VPWR VPWR U$$978/A sky130_fd_sc_hd__a22o_1
XU$$1127 U$$1127/A U$$1163/B VGND VGND VPWR VPWR U$$1127/X sky130_fd_sc_hd__xor2_1
XU$$988 U$$988/A U$$990/B VGND VGND VPWR VPWR U$$988/X sky130_fd_sc_hd__xor2_1
XU$$999 U$$999/A1 U$$999/A2 U$$999/B1 U$$999/B2 VGND VGND VPWR VPWR U$$999/X sky130_fd_sc_hd__a22o_1
XU$$1138 U$$42/A1 U$$1174/A2 U$$44/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1139/A sky130_fd_sc_hd__a22o_1
XFILLER_71_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1149 U$$1149/A U$$1171/B VGND VGND VPWR VPWR U$$1149/X sky130_fd_sc_hd__xor2_1
XFILLER_43_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1250 U$$651/B VGND VGND VPWR VPWR U$$684/A sky130_fd_sc_hd__buf_6
Xfanout1261 U$$4294/B VGND VGND VPWR VPWR U$$4292/B sky130_fd_sc_hd__buf_6
XFILLER_22_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_2_29_3 U$$1262/X U$$1395/X VGND VGND VPWR VPWR dadda_fa_3_30_2/B dadda_fa_4_29_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1272 fanout1279/X VGND VGND VPWR VPWR U$$4175/B sky130_fd_sc_hd__buf_6
XFILLER_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1283 U$$410/A VGND VGND VPWR VPWR U$$407/B sky130_fd_sc_hd__clkbuf_8
XFILLER_93_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1294 U$$4058/B VGND VGND VPWR VPWR U$$4098/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_42_3 input193/X dadda_fa_2_42_3/B dadda_fa_2_42_3/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_43_1/B dadda_fa_3_42_3/B sky130_fd_sc_hd__fa_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3030 U$$3030/A1 U$$3066/A2 U$$3030/B1 U$$3066/B2 VGND VGND VPWR VPWR U$$3031/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3041 U$$3041/A U$$3077/B VGND VGND VPWR VPWR U$$3041/X sky130_fd_sc_hd__xor2_1
XU$$3052 U$$3189/A1 U$$3072/A2 U$$999/A1 U$$3072/B2 VGND VGND VPWR VPWR U$$3053/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3063 U$$3063/A U$$3107/B VGND VGND VPWR VPWR U$$3063/X sky130_fd_sc_hd__xor2_1
XFILLER_53_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_35_2 U$$1141/X U$$1274/X U$$1407/X VGND VGND VPWR VPWR dadda_fa_3_36_1/A
+ dadda_fa_3_35_3/A sky130_fd_sc_hd__fa_1
XU$$3074 U$$745/A1 U$$3124/A2 U$$745/B1 U$$3124/B2 VGND VGND VPWR VPWR U$$3075/A sky130_fd_sc_hd__a22o_1
XU$$2340 U$$2340/A U$$2416/B VGND VGND VPWR VPWR U$$2340/X sky130_fd_sc_hd__xor2_1
XU$$3085 U$$3085/A U$$3150/A VGND VGND VPWR VPWR U$$3085/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_12_1 dadda_fa_5_12_1/A dadda_fa_5_12_1/B dadda_ha_4_12_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_13_0/B dadda_fa_7_12_0/A sky130_fd_sc_hd__fa_1
XU$$2351 U$$2625/A1 U$$2395/A2 U$$983/A1 U$$2395/B2 VGND VGND VPWR VPWR U$$2352/A
+ sky130_fd_sc_hd__a22o_1
XU$$3096 U$$3370/A1 U$$3108/A2 U$$3370/B1 U$$3108/B2 VGND VGND VPWR VPWR U$$3097/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_28_1 U$$462/X U$$595/X U$$728/X VGND VGND VPWR VPWR dadda_fa_3_29_2/A
+ dadda_fa_3_28_3/B sky130_fd_sc_hd__fa_1
XU$$2362 U$$2362/A U$$2396/B VGND VGND VPWR VPWR U$$2362/X sky130_fd_sc_hd__xor2_1
XU$$2373 U$$2647/A1 U$$2413/A2 U$$183/A1 U$$2413/B2 VGND VGND VPWR VPWR U$$2374/A
+ sky130_fd_sc_hd__a22o_1
XU$$2384 U$$2384/A U$$2412/B VGND VGND VPWR VPWR U$$2384/X sky130_fd_sc_hd__xor2_1
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1650 U$$1650/A1 U$$1698/A2 U$$2748/A1 U$$1698/B2 VGND VGND VPWR VPWR U$$1651/A
+ sky130_fd_sc_hd__a22o_1
XU$$2395 U$$3628/A1 U$$2395/A2 U$$3628/B1 U$$2395/B2 VGND VGND VPWR VPWR U$$2396/A
+ sky130_fd_sc_hd__a22o_1
XU$$1661 U$$1661/A U$$1697/B VGND VGND VPWR VPWR U$$1661/X sky130_fd_sc_hd__xor2_1
XU$$1672 U$$28/A1 U$$1702/A2 U$$30/A1 U$$1702/B2 VGND VGND VPWR VPWR U$$1673/A sky130_fd_sc_hd__a22o_1
XU$$1683 U$$1683/A U$$1699/B VGND VGND VPWR VPWR U$$1683/X sky130_fd_sc_hd__xor2_1
XU$$1694 U$$596/B1 U$$1696/A2 U$$598/B1 U$$1696/B2 VGND VGND VPWR VPWR U$$1695/A sky130_fd_sc_hd__a22o_1
XFILLER_147_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$302 final_adder.U$$304/B final_adder.U$$302/B VGND VGND VPWR VPWR
+ final_adder.U$$428/B sky130_fd_sc_hd__and2_1
XFILLER_58_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$313 final_adder.U$$312/B final_adder.U$$187/X final_adder.U$$185/X
+ VGND VGND VPWR VPWR final_adder.U$$313/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$324 final_adder.U$$326/B final_adder.U$$324/B VGND VGND VPWR VPWR
+ final_adder.U$$450/B sky130_fd_sc_hd__and2_1
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$335 final_adder.U$$334/B final_adder.U$$209/X final_adder.U$$207/X
+ VGND VGND VPWR VPWR final_adder.U$$335/X sky130_fd_sc_hd__a21o_1
XFILLER_29_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$346 final_adder.U$$348/B final_adder.U$$346/B VGND VGND VPWR VPWR
+ final_adder.U$$472/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$357 final_adder.U$$356/B final_adder.U$$231/X final_adder.U$$229/X
+ VGND VGND VPWR VPWR final_adder.U$$357/X sky130_fd_sc_hd__a21o_1
XFILLER_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$368 final_adder.U$$370/B final_adder.U$$368/B VGND VGND VPWR VPWR
+ final_adder.U$$494/B sky130_fd_sc_hd__and2_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$207 U$$481/A1 U$$207/A2 U$$72/A1 U$$207/B2 VGND VGND VPWR VPWR U$$208/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$379 final_adder.U$$378/B final_adder.U$$253/X final_adder.U$$251/X
+ VGND VGND VPWR VPWR final_adder.U$$379/X sky130_fd_sc_hd__a21o_1
XU$$218 U$$218/A U$$220/B VGND VGND VPWR VPWR U$$218/X sky130_fd_sc_hd__xor2_1
XFILLER_84_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$229 U$$92/A1 U$$229/A2 U$$94/A1 U$$229/B2 VGND VGND VPWR VPWR U$$230/A sky130_fd_sc_hd__a22o_1
XFILLER_55_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_111_0 U$$3287/Y U$$3421/X U$$3554/X VGND VGND VPWR VPWR dadda_fa_4_112_1/A
+ dadda_fa_4_111_2/A sky130_fd_sc_hd__fa_1
XFILLER_5_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_52_2 dadda_fa_3_52_2/A dadda_fa_3_52_2/B dadda_fa_3_52_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_1/A dadda_fa_4_52_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_0_68_2 U$$1074/X U$$1207/X U$$1340/X VGND VGND VPWR VPWR dadda_fa_1_69_6/B
+ dadda_fa_1_68_8/A sky130_fd_sc_hd__fa_1
XFILLER_76_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_45_1 dadda_fa_3_45_1/A dadda_fa_3_45_1/B dadda_fa_3_45_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_0/CIN dadda_fa_4_45_2/A sky130_fd_sc_hd__fa_1
XFILLER_76_776 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_22_0 dadda_fa_6_22_0/A dadda_fa_6_22_0/B dadda_fa_6_22_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_23_0/B dadda_fa_7_22_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_38_0 dadda_fa_3_38_0/A dadda_fa_3_38_0/B dadda_fa_3_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_0/B dadda_fa_4_38_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$891 final_adder.U$$794/X final_adder.U$$503/X final_adder.U$$795/X
+ VGND VGND VPWR VPWR final_adder.U$$891/X sky130_fd_sc_hd__a21o_1
XU$$730 U$$730/A U$$764/B VGND VGND VPWR VPWR U$$730/X sky130_fd_sc_hd__xor2_1
XU$$741 U$$741/A1 U$$743/A2 U$$880/A1 U$$743/B2 VGND VGND VPWR VPWR U$$742/A sky130_fd_sc_hd__a22o_1
XU$$752 U$$752/A U$$768/B VGND VGND VPWR VPWR U$$752/X sky130_fd_sc_hd__xor2_1
XU$$763 U$$900/A1 U$$763/A2 U$$900/B1 U$$763/B2 VGND VGND VPWR VPWR U$$764/A sky130_fd_sc_hd__a22o_1
XU$$774 U$$774/A U$$774/B VGND VGND VPWR VPWR U$$774/X sky130_fd_sc_hd__xor2_1
XU$$785 U$$920/B1 U$$817/A2 U$$787/A1 U$$817/B2 VGND VGND VPWR VPWR U$$786/A sky130_fd_sc_hd__a22o_1
XFILLER_32_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$796 U$$796/A U$$804/B VGND VGND VPWR VPWR U$$796/X sky130_fd_sc_hd__xor2_1
XFILLER_72_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_97_4 U$$3925/X U$$4058/X U$$4191/X VGND VGND VPWR VPWR dadda_fa_3_98_1/CIN
+ dadda_fa_3_97_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout509 U$$3257/A2 VGND VGND VPWR VPWR U$$3251/A2 sky130_fd_sc_hd__buf_2
XFILLER_99_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1080 input83/X VGND VGND VPWR VPWR U$$3072/B1 sky130_fd_sc_hd__buf_4
Xfanout1091 U$$4442/A1 VGND VGND VPWR VPWR U$$4440/B1 sky130_fd_sc_hd__buf_4
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_40_0 U$$1550/X U$$1683/X U$$1816/X VGND VGND VPWR VPWR dadda_fa_3_41_0/B
+ dadda_fa_3_40_2/B sky130_fd_sc_hd__fa_1
XFILLER_54_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2170 U$$2170/A U$$2192/A VGND VGND VPWR VPWR U$$2170/X sky130_fd_sc_hd__xor2_1
XFILLER_50_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2181 U$$4508/B1 U$$2181/A2 U$$4375/A1 U$$2181/B2 VGND VGND VPWR VPWR U$$2182/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2192 U$$2192/A VGND VGND VPWR VPWR U$$2192/Y sky130_fd_sc_hd__inv_1
XFILLER_22_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1480 U$$521/A1 U$$1480/A2 U$$521/B1 U$$1480/B2 VGND VGND VPWR VPWR U$$1481/A sky130_fd_sc_hd__a22o_1
XFILLER_50_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$1491 U$$1491/A U$$1491/B VGND VGND VPWR VPWR U$$1491/X sky130_fd_sc_hd__xor2_1
XFILLER_22_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_85_2 U$$2305/X U$$2438/X U$$2571/X VGND VGND VPWR VPWR dadda_fa_2_86_3/A
+ dadda_fa_2_85_5/A sky130_fd_sc_hd__fa_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$417_1833 VGND VGND VPWR VPWR U$$417_1833/HI U$$417/A1 sky130_fd_sc_hd__conb_1
Xdadda_fa_4_62_1 dadda_fa_4_62_1/A dadda_fa_4_62_1/B dadda_fa_4_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_63_0/B dadda_fa_5_62_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_78_1 U$$1626/X U$$1759/X U$$1892/X VGND VGND VPWR VPWR dadda_fa_2_79_0/CIN
+ dadda_fa_2_78_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_77_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_55_0 dadda_fa_4_55_0/A dadda_fa_4_55_0/B dadda_fa_4_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_56_0/A dadda_fa_5_55_1/A sky130_fd_sc_hd__fa_1
XFILLER_103_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$110 _406_/Q _278_/Q VGND VGND VPWR VPWR final_adder.U$$915/B1 final_adder.U$$144/A
+ sky130_fd_sc_hd__ha_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$121 _417_/Q _289_/Q VGND VGND VPWR VPWR final_adder.U$$135/B1 final_adder.U$$134/B
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$132 final_adder.U$$132/A final_adder.U$$132/B VGND VGND VPWR VPWR
+ final_adder.U$$260/B sky130_fd_sc_hd__and2_1
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$143 final_adder.U$$142/B final_adder.U$$913/B1 final_adder.U$$143/B1
+ VGND VGND VPWR VPWR final_adder.U$$143/X sky130_fd_sc_hd__a21o_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$154 final_adder.U$$154/A final_adder.U$$154/B VGND VGND VPWR VPWR
+ final_adder.U$$282/B sky130_fd_sc_hd__and2_1
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$165 final_adder.U$$164/B final_adder.U$$935/B1 final_adder.U$$165/B1
+ VGND VGND VPWR VPWR final_adder.U$$165/X sky130_fd_sc_hd__a21o_1
XFILLER_46_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$176 final_adder.U$$176/A final_adder.U$$176/B VGND VGND VPWR VPWR
+ final_adder.U$$304/B sky130_fd_sc_hd__and2_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$187 final_adder.U$$186/B final_adder.U$$957/B1 final_adder.U$$187/B1
+ VGND VGND VPWR VPWR final_adder.U$$187/X sky130_fd_sc_hd__a21o_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$198 final_adder.U$$198/A final_adder.U$$198/B VGND VGND VPWR VPWR
+ final_adder.U$$326/B sky130_fd_sc_hd__and2_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_382_ _382_/CLK _382_/D VGND VGND VPWR VPWR _382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_0_74_2 U$$1485/X U$$1618/X VGND VGND VPWR VPWR dadda_fa_1_75_8/B dadda_fa_2_74_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_73_0 U$$684/Y U$$818/X U$$951/X VGND VGND VPWR VPWR dadda_fa_1_74_7/B
+ dadda_fa_1_73_8/B sky130_fd_sc_hd__fa_1
XFILLER_110_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput150 c[119] VGND VGND VPWR VPWR input150/X sky130_fd_sc_hd__buf_2
Xinput161 c[13] VGND VGND VPWR VPWR input161/X sky130_fd_sc_hd__clkbuf_4
Xinput172 c[23] VGND VGND VPWR VPWR input172/X sky130_fd_sc_hd__buf_2
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput183 c[33] VGND VGND VPWR VPWR input183/X sky130_fd_sc_hd__buf_2
Xinput194 c[43] VGND VGND VPWR VPWR input194/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$560 U$$697/A1 U$$610/A2 U$$14/A1 U$$610/B2 VGND VGND VPWR VPWR U$$561/A sky130_fd_sc_hd__a22o_1
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$571 U$$571/A U$$639/B VGND VGND VPWR VPWR U$$571/X sky130_fd_sc_hd__xor2_1
XU$$582 U$$34/A1 U$$638/A2 U$$36/A1 U$$638/B2 VGND VGND VPWR VPWR U$$583/A sky130_fd_sc_hd__a22o_1
XFILLER_17_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$593 U$$593/A U$$631/B VGND VGND VPWR VPWR U$$593/X sky130_fd_sc_hd__xor2_1
XFILLER_60_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_95_1 U$$2990/X U$$3123/X U$$3256/X VGND VGND VPWR VPWR dadda_fa_3_96_0/CIN
+ dadda_fa_3_95_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_133_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_72_0 dadda_fa_5_72_0/A dadda_fa_5_72_0/B dadda_fa_5_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_73_0/A dadda_fa_6_72_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_88_0 U$$3508/X U$$3641/X U$$3774/X VGND VGND VPWR VPWR dadda_fa_3_89_0/B
+ dadda_fa_3_88_2/B sky130_fd_sc_hd__fa_1
XFILLER_113_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_71_8 dadda_fa_1_71_8/A dadda_fa_1_71_8/B dadda_fa_1_71_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_72_3/A dadda_fa_3_71_0/A sky130_fd_sc_hd__fa_1
XFILLER_87_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_7 dadda_fa_1_64_7/A dadda_fa_1_64_7/B dadda_fa_1_64_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_65_2/CIN dadda_fa_2_64_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_57_6 U$$3579/X U$$3712/X U$$3845/X VGND VGND VPWR VPWR dadda_fa_2_58_2/B
+ dadda_fa_2_57_5/B sky130_fd_sc_hd__fa_1
XFILLER_67_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_9_0 dadda_fa_7_9_0/A dadda_fa_7_9_0/B dadda_fa_7_9_0/CIN VGND VGND VPWR
+ VPWR _306_/D _177_/D sky130_fd_sc_hd__fa_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_87_0 dadda_fa_7_87_0/A dadda_fa_7_87_0/B dadda_fa_7_87_0/CIN VGND VGND
+ VPWR VPWR _384_/D _255_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_1_90_0 dadda_fa_1_90_0/A U$$1916/X U$$2049/X VGND VGND VPWR VPWR dadda_fa_2_91_4/A
+ dadda_fa_2_90_5/A sky130_fd_sc_hd__fa_1
XFILLER_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout840 U$$2060/X VGND VGND VPWR VPWR U$$2147/B2 sky130_fd_sc_hd__buf_6
Xfanout851 U$$2022/B2 VGND VGND VPWR VPWR U$$2052/B2 sky130_fd_sc_hd__buf_6
Xfanout862 U$$1726/B2 VGND VGND VPWR VPWR U$$1696/B2 sky130_fd_sc_hd__clkbuf_4
XU$$4308 U$$4308/A U$$4384/A VGND VGND VPWR VPWR U$$4308/X sky130_fd_sc_hd__xor2_1
Xfanout873 U$$1621/B2 VGND VGND VPWR VPWR U$$1593/B2 sky130_fd_sc_hd__buf_2
XFILLER_120_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout884 U$$213/B2 VGND VGND VPWR VPWR U$$179/B2 sky130_fd_sc_hd__clkbuf_4
XU$$4319 U$$4456/A1 U$$4325/A2 U$$4456/B1 U$$4325/B2 VGND VGND VPWR VPWR U$$4320/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout895 U$$1375/X VGND VGND VPWR VPWR U$$1480/B2 sky130_fd_sc_hd__buf_8
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3607 U$$3607/A U$$3607/B VGND VGND VPWR VPWR U$$3607/X sky130_fd_sc_hd__xor2_1
XFILLER_92_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3618 U$$3618/A1 U$$3696/A2 U$$3618/B1 U$$3696/B2 VGND VGND VPWR VPWR U$$3619/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3629 U$$3629/A U$$3641/B VGND VGND VPWR VPWR U$$3629/X sky130_fd_sc_hd__xor2_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_102_0 dadda_fa_6_102_0/A dadda_fa_6_102_0/B dadda_fa_6_102_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_103_0/B dadda_fa_7_102_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2906 U$$2906/A U$$2944/B VGND VGND VPWR VPWR U$$2906/X sky130_fd_sc_hd__xor2_1
XU$$2917 U$$999/A1 U$$2937/A2 U$$999/B1 U$$2937/B2 VGND VGND VPWR VPWR U$$2918/A sky130_fd_sc_hd__a22o_1
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2928 U$$2928/A U$$2938/B VGND VGND VPWR VPWR U$$2928/X sky130_fd_sc_hd__xor2_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2939 U$$4446/A1 U$$2977/A2 U$$4446/B1 U$$2977/B2 VGND VGND VPWR VPWR U$$2940/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_22_3 U$$1514/X U$$1570/B input171/X VGND VGND VPWR VPWR dadda_fa_4_23_1/B
+ dadda_fa_4_22_2/CIN sky130_fd_sc_hd__fa_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4407_1851 VGND VGND VPWR VPWR U$$4407_1851/HI U$$4407/B sky130_fd_sc_hd__conb_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_365_ _366_/CLK _365_/D VGND VGND VPWR VPWR _365_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_296_ _319_/CLK _296_/D VGND VGND VPWR VPWR _296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_67_5 dadda_fa_2_67_5/A dadda_fa_2_67_5/B dadda_fa_2_67_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_2/A dadda_fa_4_67_0/A sky130_fd_sc_hd__fa_1
XFILLER_96_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_930 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$390 U$$936/B1 U$$406/A2 U$$803/A1 U$$406/B2 VGND VGND VPWR VPWR U$$391/A sky130_fd_sc_hd__a22o_1
XFILLER_51_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_62_4 U$$3988/X U$$4121/X U$$4254/X VGND VGND VPWR VPWR dadda_fa_2_63_1/CIN
+ dadda_fa_2_62_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_55_3 U$$1979/X U$$2112/X U$$2245/X VGND VGND VPWR VPWR dadda_fa_2_56_1/B
+ dadda_fa_2_55_4/B sky130_fd_sc_hd__fa_1
XFILLER_170_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_32_2 dadda_fa_4_32_2/A dadda_fa_4_32_2/B dadda_fa_4_32_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_33_0/CIN dadda_fa_5_32_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_48_2 U$$901/X U$$1034/X U$$1167/X VGND VGND VPWR VPWR dadda_fa_2_49_1/CIN
+ dadda_fa_2_48_4/B sky130_fd_sc_hd__fa_1
XFILLER_55_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_25_1 dadda_fa_4_25_1/A dadda_fa_4_25_1/B dadda_fa_4_25_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_26_0/B dadda_fa_5_25_1/B sky130_fd_sc_hd__fa_1
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_18_0 U$$1107/X U$$1240/X U$$1278/B VGND VGND VPWR VPWR dadda_fa_5_19_0/A
+ dadda_fa_5_18_1/A sky130_fd_sc_hd__fa_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4437_1866 VGND VGND VPWR VPWR U$$4437_1866/HI U$$4437/B sky130_fd_sc_hd__conb_1
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1602 U$$2042/A1 VGND VGND VPWR VPWR U$$944/B1 sky130_fd_sc_hd__buf_2
XFILLER_78_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1613 U$$2860/B1 VGND VGND VPWR VPWR U$$120/B1 sky130_fd_sc_hd__buf_6
Xfanout1624 U$$4504/A1 VGND VGND VPWR VPWR U$$3817/B1 sky130_fd_sc_hd__buf_4
Xfanout1635 U$$2993/B1 VGND VGND VPWR VPWR U$$4502/A1 sky130_fd_sc_hd__buf_2
Xfanout1646 U$$388/A1 VGND VGND VPWR VPWR U$$936/A1 sky130_fd_sc_hd__buf_4
XU$$4105 U$$4240/B1 U$$4105/A2 U$$4107/A1 U$$4105/B2 VGND VGND VPWR VPWR U$$4106/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1657 U$$2578/A1 VGND VGND VPWR VPWR U$$521/B1 sky130_fd_sc_hd__buf_6
Xfanout670 U$$807/B2 VGND VGND VPWR VPWR U$$809/B2 sky130_fd_sc_hd__buf_4
XU$$4116 U$$4116/A1 U$$4158/A2 U$$4392/A1 U$$4158/B2 VGND VGND VPWR VPWR U$$4117/A
+ sky130_fd_sc_hd__a22o_1
Xfanout1668 U$$4494/A1 VGND VGND VPWR VPWR U$$4220/A1 sky130_fd_sc_hd__buf_4
XU$$4127 U$$4127/A U$$4133/B VGND VGND VPWR VPWR U$$4127/X sky130_fd_sc_hd__xor2_1
Xfanout681 U$$642/B2 VGND VGND VPWR VPWR U$$638/B2 sky130_fd_sc_hd__buf_4
Xfanout1679 fanout1680/X VGND VGND VPWR VPWR U$$4353/B1 sky130_fd_sc_hd__buf_4
XU$$4138 U$$4412/A1 U$$4244/A2 U$$4414/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4139/A
+ sky130_fd_sc_hd__a22o_1
Xfanout692 U$$4252/X VGND VGND VPWR VPWR U$$4309/B2 sky130_fd_sc_hd__buf_2
XU$$3404 U$$3815/A1 U$$3418/A2 U$$4226/B1 U$$3418/B2 VGND VGND VPWR VPWR U$$3405/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4149 U$$4149/A U$$4231/B VGND VGND VPWR VPWR U$$4149/X sky130_fd_sc_hd__xor2_1
XU$$3415 U$$3415/A U$$3417/B VGND VGND VPWR VPWR U$$3415/X sky130_fd_sc_hd__xor2_1
XU$$3426 input46/X VGND VGND VPWR VPWR U$$3428/B sky130_fd_sc_hd__inv_1
XFILLER_92_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3437 U$$971/A1 U$$3439/A2 U$$562/A1 U$$3439/B2 VGND VGND VPWR VPWR U$$3438/A sky130_fd_sc_hd__a22o_1
XFILLER_37_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2703 U$$2840/A1 U$$2707/A2 U$$2840/B1 U$$2707/B2 VGND VGND VPWR VPWR U$$2704/A
+ sky130_fd_sc_hd__a22o_1
XU$$3448 U$$3448/A U$$3482/B VGND VGND VPWR VPWR U$$3448/X sky130_fd_sc_hd__xor2_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2714 U$$2714/A U$$2739/A VGND VGND VPWR VPWR U$$2714/X sky130_fd_sc_hd__xor2_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3459 U$$3870/A1 U$$3471/A2 U$$3870/B1 U$$3471/B2 VGND VGND VPWR VPWR U$$3460/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2725 U$$120/B1 U$$2737/A2 U$$946/A1 U$$2737/B2 VGND VGND VPWR VPWR U$$2726/A sky130_fd_sc_hd__a22o_1
XU$$2736 U$$2736/A U$$2738/B VGND VGND VPWR VPWR U$$2736/X sky130_fd_sc_hd__xor2_1
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2747 U$$2747/A U$$2805/B VGND VGND VPWR VPWR U$$2747/X sky130_fd_sc_hd__xor2_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2758 U$$2758/A1 U$$2798/A2 U$$2758/B1 U$$2798/B2 VGND VGND VPWR VPWR U$$2759/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_0 U$$47/X U$$180/X U$$313/X VGND VGND VPWR VPWR dadda_fa_4_21_0/B dadda_fa_4_20_1/CIN
+ sky130_fd_sc_hd__fa_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2769 U$$2769/A U$$2811/B VGND VGND VPWR VPWR U$$2769/X sky130_fd_sc_hd__xor2_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_417_ _420_/CLK _417_/D VGND VGND VPWR VPWR _417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_348_ _348_/CLK _348_/D VGND VGND VPWR VPWR _348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_999 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_279_ _408_/CLK _279_/D VGND VGND VPWR VPWR _279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1000 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_72_3 dadda_fa_2_72_3/A dadda_fa_2_72_3/B dadda_fa_2_72_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_1/B dadda_fa_3_72_3/B sky130_fd_sc_hd__fa_1
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_65_2 dadda_fa_2_65_2/A dadda_fa_2_65_2/B dadda_fa_2_65_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_1/A dadda_fa_3_65_3/A sky130_fd_sc_hd__fa_1
XFILLER_68_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$709 final_adder.U$$708/B final_adder.U$$605/X final_adder.U$$589/X
+ VGND VGND VPWR VPWR final_adder.U$$709/X sky130_fd_sc_hd__a21o_1
XFILLER_69_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_42_1 dadda_fa_5_42_1/A dadda_fa_5_42_1/B dadda_fa_5_42_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_43_0/B dadda_fa_7_42_0/A sky130_fd_sc_hd__fa_2
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_58_1 dadda_fa_2_58_1/A dadda_fa_2_58_1/B dadda_fa_2_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_0/CIN dadda_fa_3_58_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_65_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_35_0 dadda_fa_5_35_0/A dadda_fa_5_35_0/B dadda_fa_5_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_36_0/A dadda_fa_6_35_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_37_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3960 U$$3960/A1 U$$3960/A2 U$$3960/B1 U$$3960/B2 VGND VGND VPWR VPWR U$$3961/A
+ sky130_fd_sc_hd__a22o_1
XU$$3971 U$$3971/A U$$3972/A VGND VGND VPWR VPWR U$$3971/X sky130_fd_sc_hd__xor2_1
XU$$3982 U$$3982/A U$$4006/B VGND VGND VPWR VPWR U$$3982/X sky130_fd_sc_hd__xor2_1
XFILLER_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3993 U$$4265/B1 U$$4025/A2 U$$4132/A1 U$$4025/B2 VGND VGND VPWR VPWR U$$3994/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput262 output262/A VGND VGND VPWR VPWR o[104] sky130_fd_sc_hd__buf_2
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput273 output273/A VGND VGND VPWR VPWR o[114] sky130_fd_sc_hd__buf_2
Xoutput284 output284/A VGND VGND VPWR VPWR o[124] sky130_fd_sc_hd__buf_2
Xoutput295 output295/A VGND VGND VPWR VPWR o[19] sky130_fd_sc_hd__buf_2
XFILLER_99_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_60_1 U$$2388/X U$$2521/X U$$2654/X VGND VGND VPWR VPWR dadda_fa_2_61_0/CIN
+ dadda_fa_2_60_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_87_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_53_0 U$$379/X U$$512/X U$$645/X VGND VGND VPWR VPWR dadda_fa_2_54_0/B
+ dadda_fa_2_53_3/B sky130_fd_sc_hd__fa_1
XFILLER_83_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1309 U$$76/A1 U$$1309/A2 U$$78/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1310/A sky130_fd_sc_hd__a22o_1
XFILLER_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_202_ _344_/CLK _202_/D VGND VGND VPWR VPWR _202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1103 final_adder.U$$176/B final_adder.U$$947/X VGND VGND VPWR VPWR
+ output361/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1114 final_adder.U$$164/A final_adder.U$$873/X VGND VGND VPWR VPWR
+ output374/A sky130_fd_sc_hd__xor2_1
XFILLER_11_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1125 final_adder.U$$154/B final_adder.U$$925/X VGND VGND VPWR VPWR
+ output259/A sky130_fd_sc_hd__xor2_1
XFILLER_137_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1136 final_adder.U$$142/A final_adder.U$$851/X VGND VGND VPWR VPWR
+ output271/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1147 final_adder.U$$132/B final_adder.U$$903/X VGND VGND VPWR VPWR
+ output283/A sky130_fd_sc_hd__xor2_1
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_82_2 dadda_fa_3_82_2/A dadda_fa_3_82_2/B dadda_fa_3_82_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_1/A dadda_fa_4_82_2/B sky130_fd_sc_hd__fa_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_75_1 dadda_fa_3_75_1/A dadda_fa_3_75_1/B dadda_fa_3_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_0/CIN dadda_fa_4_75_2/A sky130_fd_sc_hd__fa_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_52_0 dadda_fa_6_52_0/A dadda_fa_6_52_0/B dadda_fa_6_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_53_0/B dadda_fa_7_52_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_68_0 dadda_fa_3_68_0/A dadda_fa_3_68_0/B dadda_fa_3_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_0/B dadda_fa_4_68_1/CIN sky130_fd_sc_hd__fa_1
Xfanout1410 input33/X VGND VGND VPWR VPWR U$$2745/A2 sky130_fd_sc_hd__buf_6
Xfanout1421 U$$821/A VGND VGND VPWR VPWR U$$768/B sky130_fd_sc_hd__buf_6
Xfanout1432 U$$2408/B VGND VGND VPWR VPWR U$$2446/B sky130_fd_sc_hd__buf_4
XFILLER_66_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1443 U$$2273/B VGND VGND VPWR VPWR U$$2283/B sky130_fd_sc_hd__buf_4
Xfanout1454 U$$2168/B VGND VGND VPWR VPWR U$$2192/A sky130_fd_sc_hd__buf_4
XU$$2335_1802 VGND VGND VPWR VPWR U$$2335_1802/HI U$$2335/A1 sky130_fd_sc_hd__conb_1
Xfanout1465 U$$2054/A VGND VGND VPWR VPWR U$$2031/B sky130_fd_sc_hd__buf_6
Xfanout1476 input20/X VGND VGND VPWR VPWR U$$1916/B sky130_fd_sc_hd__buf_6
XFILLER_47_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1487 U$$1594/B VGND VGND VPWR VPWR U$$1568/B sky130_fd_sc_hd__buf_4
Xfanout1498 U$$1455/B VGND VGND VPWR VPWR U$$1461/B sky130_fd_sc_hd__buf_6
XU$$3201 U$$4295/B1 U$$3207/A2 U$$4162/A1 U$$3207/B2 VGND VGND VPWR VPWR U$$3202/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3212 U$$3212/A U$$3258/B VGND VGND VPWR VPWR U$$3212/X sky130_fd_sc_hd__xor2_1
XU$$3223 U$$3495/B1 U$$3241/A2 U$$3499/A1 U$$3241/B2 VGND VGND VPWR VPWR U$$3224/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_111_2 dadda_fa_4_111_2/A dadda_fa_4_111_2/B dadda_fa_4_111_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_112_0/CIN dadda_fa_5_111_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_93_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$16 _312_/Q _184_/Q VGND VGND VPWR VPWR final_adder.U$$239/A2 final_adder.U$$238/A
+ sky130_fd_sc_hd__ha_1
XU$$3234 U$$3234/A U$$3242/B VGND VGND VPWR VPWR U$$3234/X sky130_fd_sc_hd__xor2_1
XU$$3245 U$$3382/A1 U$$3245/A2 U$$3382/B1 U$$3245/B2 VGND VGND VPWR VPWR U$$3246/A
+ sky130_fd_sc_hd__a22o_1
XU$$2500 U$$3048/A1 U$$2546/A2 U$$3048/B1 U$$2546/B2 VGND VGND VPWR VPWR U$$2501/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$27 _323_/Q _195_/Q VGND VGND VPWR VPWR final_adder.U$$229/B1 final_adder.U$$228/B
+ sky130_fd_sc_hd__ha_1
XU$$2511 U$$2511/A U$$2549/B VGND VGND VPWR VPWR U$$2511/X sky130_fd_sc_hd__xor2_1
XU$$3256 U$$3256/A U$$3258/B VGND VGND VPWR VPWR U$$3256/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$38 _334_/Q _206_/Q VGND VGND VPWR VPWR final_adder.U$$987/B1 final_adder.U$$216/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_4_104_1 dadda_fa_4_104_1/A dadda_fa_4_104_1/B dadda_fa_4_104_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_105_0/B dadda_fa_5_104_1/B sky130_fd_sc_hd__fa_1
XU$$3267 U$$3815/A1 U$$3285/A2 U$$3817/A1 U$$3285/B2 VGND VGND VPWR VPWR U$$3268/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2522 U$$3205/B1 U$$2532/A2 U$$3072/A1 U$$2532/B2 VGND VGND VPWR VPWR U$$2523/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$49 _345_/Q _217_/Q VGND VGND VPWR VPWR final_adder.U$$207/B1 final_adder.U$$206/B
+ sky130_fd_sc_hd__ha_1
XU$$2533 U$$2533/A U$$2541/B VGND VGND VPWR VPWR U$$2533/X sky130_fd_sc_hd__xor2_1
XFILLER_62_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3278 U$$3278/A U$$3286/B VGND VGND VPWR VPWR U$$3278/X sky130_fd_sc_hd__xor2_1
XU$$3289 input43/X VGND VGND VPWR VPWR U$$3291/B sky130_fd_sc_hd__inv_1
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2544 U$$4462/A1 U$$2546/A2 U$$3916/A1 U$$2546/B2 VGND VGND VPWR VPWR U$$2545/A
+ sky130_fd_sc_hd__a22o_1
XU$$1810 U$$1810/A U$$1836/B VGND VGND VPWR VPWR U$$1810/X sky130_fd_sc_hd__xor2_1
XU$$2555 U$$2555/A U$$2591/B VGND VGND VPWR VPWR U$$2555/X sky130_fd_sc_hd__xor2_1
XU$$2566 U$$2840/A1 U$$2574/A2 U$$2840/B1 U$$2574/B2 VGND VGND VPWR VPWR U$$2567/A
+ sky130_fd_sc_hd__a22o_1
XU$$1821 U$$997/B1 U$$1829/A2 U$$864/A1 U$$1829/B2 VGND VGND VPWR VPWR U$$1822/A sky130_fd_sc_hd__a22o_1
XU$$1832 U$$1832/A U$$1832/B VGND VGND VPWR VPWR U$$1832/X sky130_fd_sc_hd__xor2_1
XU$$2577 U$$2577/A U$$2603/A VGND VGND VPWR VPWR U$$2577/X sky130_fd_sc_hd__xor2_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2588 U$$3684/A1 U$$2600/A2 U$$3684/B1 U$$2600/B2 VGND VGND VPWR VPWR U$$2589/A
+ sky130_fd_sc_hd__a22o_1
XU$$1843 U$$745/B1 U$$1881/A2 U$$612/A1 U$$1881/B2 VGND VGND VPWR VPWR U$$1844/A sky130_fd_sc_hd__a22o_1
XU$$1854 U$$1854/A U$$1854/B VGND VGND VPWR VPWR U$$1854/X sky130_fd_sc_hd__xor2_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2599 U$$2599/A U$$2602/A VGND VGND VPWR VPWR U$$2599/X sky130_fd_sc_hd__xor2_1
XU$$1865 U$$3370/B1 U$$1909/A2 U$$3372/B1 U$$1909/B2 VGND VGND VPWR VPWR U$$1866/A
+ sky130_fd_sc_hd__a22o_1
XU$$1876 U$$1876/A U$$1916/B VGND VGND VPWR VPWR U$$1876/X sky130_fd_sc_hd__xor2_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1887 U$$4353/A1 U$$1915/A2 U$$4353/B1 U$$1915/B2 VGND VGND VPWR VPWR U$$1888/A
+ sky130_fd_sc_hd__a22o_1
XU$$1898 U$$1898/A U$$1910/B VGND VGND VPWR VPWR U$$1898/X sky130_fd_sc_hd__xor2_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_125_0 dadda_fa_7_125_0/A dadda_fa_7_125_0/B dadda_fa_7_125_0/CIN VGND
+ VGND VPWR VPWR _422_/D _293_/D sky130_fd_sc_hd__fa_1
XFILLER_174_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_70_0 dadda_fa_2_70_0/A dadda_fa_2_70_0/B dadda_fa_2_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_0/B dadda_fa_3_70_2/B sky130_fd_sc_hd__fa_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$517 final_adder.U$$516/B final_adder.U$$401/X final_adder.U$$393/X
+ VGND VGND VPWR VPWR final_adder.U$$517/X sky130_fd_sc_hd__a21o_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$528 final_adder.U$$536/B final_adder.U$$528/B VGND VGND VPWR VPWR
+ final_adder.U$$648/B sky130_fd_sc_hd__and2_1
XFILLER_69_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$539 final_adder.U$$538/B final_adder.U$$423/X final_adder.U$$415/X
+ VGND VGND VPWR VPWR final_adder.U$$539/X sky130_fd_sc_hd__a21o_1
XFILLER_72_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4480 U$$4480/A1 U$$4388/X U$$4482/A1 U$$4488/B2 VGND VGND VPWR VPWR U$$4481/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4491 U$$4491/A U$$4491/B VGND VGND VPWR VPWR U$$4491/X sky130_fd_sc_hd__xor2_1
XFILLER_80_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3790 U$$3790/A U$$3790/B VGND VGND VPWR VPWR U$$3790/X sky130_fd_sc_hd__xor2_1
XFILLER_80_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2874_1811 VGND VGND VPWR VPWR U$$2874_1811/HI U$$2874/B1 sky130_fd_sc_hd__conb_1
Xdadda_fa_4_92_1 dadda_fa_4_92_1/A dadda_fa_4_92_1/B dadda_fa_4_92_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_93_0/B dadda_fa_5_92_1/B sky130_fd_sc_hd__fa_1
XFILLER_109_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_85_0 dadda_fa_4_85_0/A dadda_fa_4_85_0/B dadda_fa_4_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_86_0/A dadda_fa_5_85_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_106_3 dadda_fa_3_106_3/A dadda_fa_3_106_3/B dadda_fa_3_106_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_107_1/B dadda_fa_4_106_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_107_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$901 U$$901/A U$$925/B VGND VGND VPWR VPWR U$$901/X sky130_fd_sc_hd__xor2_1
XU$$912 U$$912/A1 U$$952/A2 U$$914/A1 U$$952/B2 VGND VGND VPWR VPWR U$$913/A sky130_fd_sc_hd__a22o_1
XU$$923 U$$923/A U$$943/B VGND VGND VPWR VPWR U$$923/X sky130_fd_sc_hd__xor2_1
XFILLER_28_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$934 U$$934/A1 U$$942/A2 U$$936/A1 U$$942/B2 VGND VGND VPWR VPWR U$$935/A sky130_fd_sc_hd__a22o_1
XU$$945 U$$945/A U$$958/A VGND VGND VPWR VPWR U$$945/X sky130_fd_sc_hd__xor2_1
XU$$956 U$$956/A1 U$$956/A2 U$$956/B1 U$$956/B2 VGND VGND VPWR VPWR U$$957/A sky130_fd_sc_hd__a22o_1
XU$$1106 U$$969/A1 U$$1174/A2 U$$971/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1107/A sky130_fd_sc_hd__a22o_1
XU$$967 U$$967/A1 U$$981/A2 U$$969/A1 U$$981/B2 VGND VGND VPWR VPWR U$$968/A sky130_fd_sc_hd__a22o_1
XU$$1117 U$$1117/A U$$1171/B VGND VGND VPWR VPWR U$$1117/X sky130_fd_sc_hd__xor2_1
XU$$978 U$$978/A U$$980/B VGND VGND VPWR VPWR U$$978/X sky130_fd_sc_hd__xor2_1
XU$$1128 U$$991/A1 U$$1164/A2 U$$993/A1 U$$1164/B2 VGND VGND VPWR VPWR U$$1129/A sky130_fd_sc_hd__a22o_1
XU$$989 U$$989/A1 U$$999/A2 U$$989/B1 U$$999/B2 VGND VGND VPWR VPWR U$$990/A sky130_fd_sc_hd__a22o_1
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1139 U$$1139/A U$$1175/B VGND VGND VPWR VPWR U$$1139/X sky130_fd_sc_hd__xor2_1
XFILLER_71_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_914 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1240 U$$3979/B1 VGND VGND VPWR VPWR U$$828/B1 sky130_fd_sc_hd__clkbuf_2
Xfanout1251 input64/X VGND VGND VPWR VPWR U$$651/B sky130_fd_sc_hd__buf_8
Xfanout1262 input60/X VGND VGND VPWR VPWR U$$4294/B sky130_fd_sc_hd__buf_4
Xfanout1273 fanout1279/X VGND VGND VPWR VPWR U$$4247/A sky130_fd_sc_hd__buf_4
Xfanout1284 input56/X VGND VGND VPWR VPWR U$$410/A sky130_fd_sc_hd__buf_6
XU$$4489_1892 VGND VGND VPWR VPWR U$$4489_1892/HI U$$4489/B sky130_fd_sc_hd__conb_1
Xfanout1295 fanout1299/X VGND VGND VPWR VPWR U$$4108/B sky130_fd_sc_hd__buf_2
XFILLER_93_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_42_4 dadda_fa_2_42_4/A dadda_fa_2_42_4/B dadda_fa_2_42_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_43_1/CIN dadda_fa_3_42_3/CIN sky130_fd_sc_hd__fa_1
XU$$3020 U$$3020/A1 U$$3066/A2 U$$3022/A1 U$$3066/B2 VGND VGND VPWR VPWR U$$3021/A
+ sky130_fd_sc_hd__a22o_1
XU$$3031 U$$3031/A U$$3073/B VGND VGND VPWR VPWR U$$3031/X sky130_fd_sc_hd__xor2_1
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3042 U$$4412/A1 U$$3122/A2 U$$4414/A1 U$$3122/B2 VGND VGND VPWR VPWR U$$3043/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3053 U$$3053/A U$$3073/B VGND VGND VPWR VPWR U$$3053/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_35_3 U$$1540/X U$$1673/X U$$1806/X VGND VGND VPWR VPWR dadda_fa_3_36_1/B
+ dadda_fa_3_35_3/B sky130_fd_sc_hd__fa_1
XU$$3064 U$$4295/B1 U$$3072/A2 U$$4162/A1 U$$3072/B2 VGND VGND VPWR VPWR U$$3065/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2330 input28/X VGND VGND VPWR VPWR U$$2332/B sky130_fd_sc_hd__inv_1
XU$$3075 U$$3075/A U$$3077/B VGND VGND VPWR VPWR U$$3075/X sky130_fd_sc_hd__xor2_1
XFILLER_90_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2341 U$$971/A1 U$$2415/A2 U$$973/A1 U$$2415/B2 VGND VGND VPWR VPWR U$$2342/A sky130_fd_sc_hd__a22o_1
XU$$3086 U$$4456/A1 U$$3148/A2 U$$4456/B1 U$$3148/B2 VGND VGND VPWR VPWR U$$3087/A
+ sky130_fd_sc_hd__a22o_1
XU$$2352 U$$2352/A U$$2396/B VGND VGND VPWR VPWR U$$2352/X sky130_fd_sc_hd__xor2_1
XU$$3097 U$$3097/A U$$3107/B VGND VGND VPWR VPWR U$$3097/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_28_2 U$$861/X U$$994/X U$$1127/X VGND VGND VPWR VPWR dadda_fa_3_29_2/B
+ dadda_fa_3_28_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_90_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2363 U$$854/B1 U$$2407/A2 U$$3322/B1 U$$2407/B2 VGND VGND VPWR VPWR U$$2364/A
+ sky130_fd_sc_hd__a22o_1
XU$$2374 U$$2374/A U$$2416/B VGND VGND VPWR VPWR U$$2374/X sky130_fd_sc_hd__xor2_1
XU$$1640 U$$1640/A U$$1644/A VGND VGND VPWR VPWR U$$1640/X sky130_fd_sc_hd__xor2_1
XU$$2385 U$$3205/B1 U$$2407/A2 U$$3072/A1 U$$2407/B2 VGND VGND VPWR VPWR U$$2386/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2396 U$$2396/A U$$2396/B VGND VGND VPWR VPWR U$$2396/X sky130_fd_sc_hd__xor2_1
XU$$1651 U$$1651/A U$$1699/B VGND VGND VPWR VPWR U$$1651/X sky130_fd_sc_hd__xor2_1
XU$$1662 U$$2758/A1 U$$1698/A2 U$$2758/B1 U$$1698/B2 VGND VGND VPWR VPWR U$$1663/A
+ sky130_fd_sc_hd__a22o_1
XU$$1673 U$$1673/A U$$1703/B VGND VGND VPWR VPWR U$$1673/X sky130_fd_sc_hd__xor2_1
XU$$1684 U$$999/A1 U$$1698/A2 U$$999/B1 U$$1698/B2 VGND VGND VPWR VPWR U$$1685/A sky130_fd_sc_hd__a22o_1
XU$$1695 U$$1695/A U$$1697/B VGND VGND VPWR VPWR U$$1695/X sky130_fd_sc_hd__xor2_1
XFILLER_147_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$303 final_adder.U$$302/B final_adder.U$$177/X final_adder.U$$175/X
+ VGND VGND VPWR VPWR final_adder.U$$303/X sky130_fd_sc_hd__a21o_1
XFILLER_112_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$314 final_adder.U$$316/B final_adder.U$$314/B VGND VGND VPWR VPWR
+ final_adder.U$$440/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$325 final_adder.U$$324/B final_adder.U$$199/X final_adder.U$$197/X
+ VGND VGND VPWR VPWR final_adder.U$$325/X sky130_fd_sc_hd__a21o_1
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$336 final_adder.U$$338/B final_adder.U$$336/B VGND VGND VPWR VPWR
+ final_adder.U$$462/B sky130_fd_sc_hd__and2_1
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$347 final_adder.U$$346/B final_adder.U$$221/X final_adder.U$$219/X
+ VGND VGND VPWR VPWR final_adder.U$$347/X sky130_fd_sc_hd__a21o_1
XFILLER_29_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$358 final_adder.U$$360/B final_adder.U$$358/B VGND VGND VPWR VPWR
+ final_adder.U$$484/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$369 final_adder.U$$368/B final_adder.U$$243/X final_adder.U$$241/X
+ VGND VGND VPWR VPWR final_adder.U$$369/X sky130_fd_sc_hd__a21o_1
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$208 U$$208/A U$$210/B VGND VGND VPWR VPWR U$$208/X sky130_fd_sc_hd__xor2_1
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$219 U$$902/B1 U$$219/A2 U$$84/A1 U$$219/B2 VGND VGND VPWR VPWR U$$220/A sky130_fd_sc_hd__a22o_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_111_1 U$$3687/X U$$3820/X U$$3953/X VGND VGND VPWR VPWR dadda_fa_4_112_1/B
+ dadda_fa_4_111_2/B sky130_fd_sc_hd__fa_1
XFILLER_112_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_104_0 U$$3806/X U$$3939/X U$$4072/X VGND VGND VPWR VPWR dadda_fa_4_105_0/B
+ dadda_fa_4_104_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1028 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_999 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_52_3 dadda_fa_3_52_3/A dadda_fa_3_52_3/B dadda_fa_3_52_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_1/B dadda_fa_4_52_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_68_3 U$$1473/X U$$1606/X U$$1739/X VGND VGND VPWR VPWR dadda_fa_1_69_6/CIN
+ dadda_fa_1_68_8/B sky130_fd_sc_hd__fa_1
XFILLER_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_45_2 dadda_fa_3_45_2/A dadda_fa_3_45_2/B dadda_fa_3_45_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_1/A dadda_fa_4_45_2/B sky130_fd_sc_hd__fa_1
XFILLER_76_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$881 final_adder.U$$784/X final_adder.U$$737/X final_adder.U$$785/X
+ VGND VGND VPWR VPWR final_adder.U$$881/X sky130_fd_sc_hd__a21o_1
XU$$720 U$$720/A U$$774/B VGND VGND VPWR VPWR U$$720/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_38_1 dadda_fa_3_38_1/A dadda_fa_3_38_1/B dadda_fa_3_38_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_0/CIN dadda_fa_4_38_2/A sky130_fd_sc_hd__fa_1
XU$$731 U$$868/A1 U$$769/A2 U$$868/B1 U$$769/B2 VGND VGND VPWR VPWR U$$732/A sky130_fd_sc_hd__a22o_1
XFILLER_16_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$742 U$$742/A U$$744/B VGND VGND VPWR VPWR U$$742/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_15_0 dadda_fa_6_15_0/A dadda_fa_6_15_0/B dadda_fa_6_15_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_16_0/B dadda_fa_7_15_0/CIN sky130_fd_sc_hd__fa_1
XU$$753 U$$68/A1 U$$769/A2 U$$70/A1 U$$769/B2 VGND VGND VPWR VPWR U$$754/A sky130_fd_sc_hd__a22o_1
XU$$764 U$$764/A U$$764/B VGND VGND VPWR VPWR U$$764/X sky130_fd_sc_hd__xor2_1
XFILLER_44_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$775 U$$912/A1 U$$819/A2 U$$914/A1 U$$819/B2 VGND VGND VPWR VPWR U$$776/A sky130_fd_sc_hd__a22o_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$786 U$$786/A U$$820/B VGND VGND VPWR VPWR U$$786/X sky130_fd_sc_hd__xor2_1
XU$$797 U$$934/A1 U$$809/A2 U$$936/A1 U$$809/B2 VGND VGND VPWR VPWR U$$798/A sky130_fd_sc_hd__a22o_1
XFILLER_32_836 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_ha_3_110_3 U$$4350/X U$$4483/X VGND VGND VPWR VPWR dadda_fa_4_111_1/CIN dadda_ha_3_110_3/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_32_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_97_5 U$$4324/X U$$4457/X input253/X VGND VGND VPWR VPWR dadda_fa_3_98_2/A
+ dadda_fa_4_97_0/A sky130_fd_sc_hd__fa_1
XFILLER_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1070 U$$884/A1 VGND VGND VPWR VPWR U$$62/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1081 U$$745/A1 VGND VGND VPWR VPWR U$$882/A1 sky130_fd_sc_hd__buf_4
Xfanout1092 U$$3618/B1 VGND VGND VPWR VPWR U$$4442/A1 sky130_fd_sc_hd__buf_6
XFILLER_66_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_40_1 U$$1949/X U$$2082/X U$$2215/X VGND VGND VPWR VPWR dadda_fa_3_41_0/CIN
+ dadda_fa_3_40_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_82_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_clk _218_/CLK VGND VGND VPWR VPWR _346_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_33_0 U$$73/X U$$206/X U$$339/X VGND VGND VPWR VPWR dadda_fa_3_34_0/B dadda_fa_3_33_2/B
+ sky130_fd_sc_hd__fa_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2160 U$$2160/A U$$2168/B VGND VGND VPWR VPWR U$$2160/X sky130_fd_sc_hd__xor2_1
XU$$2171 U$$2443/B1 U$$2181/A2 U$$2310/A1 U$$2181/B2 VGND VGND VPWR VPWR U$$2172/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2182 U$$2182/A U$$2186/B VGND VGND VPWR VPWR U$$2182/X sky130_fd_sc_hd__xor2_1
XFILLER_50_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2193 input26/X VGND VGND VPWR VPWR U$$2195/B sky130_fd_sc_hd__inv_1
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1470 U$$98/B1 U$$1504/A2 U$$924/A1 U$$1504/B2 VGND VGND VPWR VPWR U$$1471/A sky130_fd_sc_hd__a22o_1
XU$$1481 U$$1481/A U$$1491/B VGND VGND VPWR VPWR U$$1481/X sky130_fd_sc_hd__xor2_1
XU$$1492 U$$944/A1 U$$1502/A2 U$$944/B1 U$$1502/B2 VGND VGND VPWR VPWR U$$1493/A sky130_fd_sc_hd__a22o_1
XFILLER_50_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_919 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_1_86_5 U$$3504/X U$$3637/X VGND VGND VPWR VPWR dadda_fa_2_87_4/B dadda_fa_3_86_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_985 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_85_3 U$$2704/X U$$2837/X U$$2970/X VGND VGND VPWR VPWR dadda_fa_2_86_3/B
+ dadda_fa_2_85_5/B sky130_fd_sc_hd__fa_1
XFILLER_131_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_62_2 dadda_fa_4_62_2/A dadda_fa_4_62_2/B dadda_fa_4_62_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_63_0/CIN dadda_fa_5_62_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_78_2 U$$2025/X U$$2158/X U$$2291/X VGND VGND VPWR VPWR dadda_fa_2_79_1/A
+ dadda_fa_2_78_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_55_1 dadda_fa_4_55_1/A dadda_fa_4_55_1/B dadda_fa_4_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_56_0/B dadda_fa_5_55_1/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$100 _396_/Q _268_/Q VGND VGND VPWR VPWR final_adder.U$$925/B1 final_adder.U$$154/A
+ sky130_fd_sc_hd__ha_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$111 _407_/Q _279_/Q VGND VGND VPWR VPWR final_adder.U$$145/B1 final_adder.U$$144/B
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_7_32_0 dadda_fa_7_32_0/A dadda_fa_7_32_0/B dadda_fa_7_32_0/CIN VGND VGND
+ VPWR VPWR _329_/D _200_/D sky130_fd_sc_hd__fa_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$122 _418_/Q _290_/Q VGND VGND VPWR VPWR final_adder.U$$903/B1 final_adder.U$$132/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_4_48_0 dadda_fa_4_48_0/A dadda_fa_4_48_0/B dadda_fa_4_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_49_0/A dadda_fa_5_48_1/A sky130_fd_sc_hd__fa_1
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$133 final_adder.U$$132/B final_adder.U$$903/B1 final_adder.U$$133/B1
+ VGND VGND VPWR VPWR final_adder.U$$133/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$144 final_adder.U$$144/A final_adder.U$$144/B VGND VGND VPWR VPWR
+ final_adder.U$$272/B sky130_fd_sc_hd__and2_1
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$155 final_adder.U$$154/B final_adder.U$$925/B1 final_adder.U$$155/B1
+ VGND VGND VPWR VPWR final_adder.U$$155/X sky130_fd_sc_hd__a21o_1
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$166 final_adder.U$$166/A final_adder.U$$166/B VGND VGND VPWR VPWR
+ final_adder.U$$294/B sky130_fd_sc_hd__and2_1
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$177 final_adder.U$$176/B final_adder.U$$947/B1 final_adder.U$$177/B1
+ VGND VGND VPWR VPWR final_adder.U$$177/X sky130_fd_sc_hd__a21o_1
XFILLER_57_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$188 final_adder.U$$188/A final_adder.U$$188/B VGND VGND VPWR VPWR
+ final_adder.U$$316/B sky130_fd_sc_hd__and2_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$199 final_adder.U$$198/B final_adder.U$$969/B1 final_adder.U$$199/B1
+ VGND VGND VPWR VPWR final_adder.U$$199/X sky130_fd_sc_hd__a21o_1
XFILLER_61_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk _388_/CLK VGND VGND VPWR VPWR _368_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_381_ _388_/CLK _381_/D VGND VGND VPWR VPWR _381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3568_1822 VGND VGND VPWR VPWR U$$3568_1822/HI U$$3568/A1 sky130_fd_sc_hd__conb_1
XFILLER_126_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_73_1 U$$1084/X U$$1217/X U$$1350/X VGND VGND VPWR VPWR dadda_fa_1_74_7/CIN
+ dadda_fa_1_73_8/CIN sky130_fd_sc_hd__fa_1
Xinput140 c[10] VGND VGND VPWR VPWR input140/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_3_50_0 dadda_fa_3_50_0/A dadda_fa_3_50_0/B dadda_fa_3_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_0/B dadda_fa_4_50_1/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_0_66_0 U$$99/B U$$272/X U$$405/X VGND VGND VPWR VPWR dadda_fa_1_67_5/B dadda_fa_1_66_7/B
+ sky130_fd_sc_hd__fa_1
Xinput151 c[11] VGND VGND VPWR VPWR input151/X sky130_fd_sc_hd__clkbuf_4
Xinput162 c[14] VGND VGND VPWR VPWR input162/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput173 c[24] VGND VGND VPWR VPWR input173/X sky130_fd_sc_hd__buf_2
Xinput184 c[34] VGND VGND VPWR VPWR input184/X sky130_fd_sc_hd__buf_2
Xinput195 c[44] VGND VGND VPWR VPWR input195/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_clk _388_/CLK VGND VGND VPWR VPWR _423_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$550 U$$669/B VGND VGND VPWR VPWR U$$550/Y sky130_fd_sc_hd__inv_1
XU$$561 U$$561/A U$$643/B VGND VGND VPWR VPWR U$$561/X sky130_fd_sc_hd__xor2_1
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$572 U$$709/A1 U$$638/A2 U$$709/B1 U$$638/B2 VGND VGND VPWR VPWR U$$573/A sky130_fd_sc_hd__a22o_1
XFILLER_32_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$583 U$$583/A U$$639/B VGND VGND VPWR VPWR U$$583/X sky130_fd_sc_hd__xor2_1
XU$$594 U$$729/B1 U$$630/A2 U$$596/A1 U$$630/B2 VGND VGND VPWR VPWR U$$595/A sky130_fd_sc_hd__a22o_1
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_95_2 U$$3389/X U$$3522/X U$$3655/X VGND VGND VPWR VPWR dadda_fa_3_96_1/A
+ dadda_fa_3_95_3/A sky130_fd_sc_hd__fa_1
XFILLER_132_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_72_1 dadda_fa_5_72_1/A dadda_fa_5_72_1/B dadda_fa_5_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_73_0/B dadda_fa_7_72_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_88_1 U$$3907/X U$$4040/X U$$4173/X VGND VGND VPWR VPWR dadda_fa_3_89_0/CIN
+ dadda_fa_3_88_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_944 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_65_0 dadda_fa_5_65_0/A dadda_fa_5_65_0/B dadda_fa_5_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_66_0/A dadda_fa_6_65_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_141_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_8 dadda_fa_1_64_8/A dadda_fa_1_64_8/B dadda_fa_1_64_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_65_3/A dadda_fa_3_64_0/A sky130_fd_sc_hd__fa_2
XFILLER_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_57_7 input209/X dadda_fa_1_57_7/B dadda_fa_1_57_7/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_58_2/CIN dadda_fa_2_57_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_19_clk _370_/CLK VGND VGND VPWR VPWR _416_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_4_0 U$$281/X U$$313/B input201/X VGND VGND VPWR VPWR dadda_fa_7_5_0/B
+ dadda_fa_7_4_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_23_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_90_1 U$$2182/X U$$2315/X U$$2448/X VGND VGND VPWR VPWR dadda_fa_2_91_4/B
+ dadda_fa_2_90_5/B sky130_fd_sc_hd__fa_1
XFILLER_105_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_83_0 U$$1369/Y U$$1503/X U$$1636/X VGND VGND VPWR VPWR dadda_fa_2_84_1/CIN
+ dadda_fa_2_83_4/A sky130_fd_sc_hd__fa_1
XFILLER_132_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout830 U$$2197/X VGND VGND VPWR VPWR U$$2272/B2 sky130_fd_sc_hd__buf_6
XU$$2472_1804 VGND VGND VPWR VPWR U$$2472_1804/HI U$$2472/A1 sky130_fd_sc_hd__conb_1
Xfanout841 U$$2181/B2 VGND VGND VPWR VPWR U$$2177/B2 sky130_fd_sc_hd__buf_6
Xfanout852 U$$1923/X VGND VGND VPWR VPWR U$$2022/B2 sky130_fd_sc_hd__buf_4
XFILLER_77_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout863 U$$1726/B2 VGND VGND VPWR VPWR U$$1698/B2 sky130_fd_sc_hd__buf_2
XU$$4309 U$$4309/A1 U$$4309/A2 U$$4446/B1 U$$4309/B2 VGND VGND VPWR VPWR U$$4310/A
+ sky130_fd_sc_hd__a22o_1
Xfanout874 U$$1587/B2 VGND VGND VPWR VPWR U$$1575/B2 sky130_fd_sc_hd__buf_4
Xfanout885 U$$207/B2 VGND VGND VPWR VPWR U$$213/B2 sky130_fd_sc_hd__buf_4
Xfanout896 U$$1327/B2 VGND VGND VPWR VPWR U$$1295/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_133_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3608 U$$4017/B1 U$$3656/A2 U$$870/A1 U$$3656/B2 VGND VGND VPWR VPWR U$$3609/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3619 U$$3619/A U$$3699/A VGND VGND VPWR VPWR U$$3619/X sky130_fd_sc_hd__xor2_1
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2907 U$$4414/A1 U$$2989/A2 U$$32/A1 U$$2989/B2 VGND VGND VPWR VPWR U$$2908/A sky130_fd_sc_hd__a22o_1
XU$$2918 U$$2918/A U$$2938/B VGND VGND VPWR VPWR U$$2918/X sky130_fd_sc_hd__xor2_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2929 U$$4162/A1 U$$2929/A2 U$$4162/B1 U$$2929/B2 VGND VGND VPWR VPWR U$$2930/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_364_ _364_/CLK _364_/D VGND VGND VPWR VPWR _364_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_295_ _388_/CLK _295_/D VGND VGND VPWR VPWR _295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_82_0 dadda_fa_6_82_0/A dadda_fa_6_82_0/B dadda_fa_6_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_83_0/B dadda_fa_7_82_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_98_0 input254/X dadda_fa_3_98_0/B dadda_fa_3_98_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_99_0/B dadda_fa_4_98_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$380 U$$517/A1 U$$386/A2 U$$517/B1 U$$386/B2 VGND VGND VPWR VPWR U$$381/A sky130_fd_sc_hd__a22o_1
XFILLER_33_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$391 U$$391/A U$$407/B VGND VGND VPWR VPWR U$$391/X sky130_fd_sc_hd__xor2_1
XFILLER_149_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_clk _201_/CLK VGND VGND VPWR VPWR _356_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_947 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_62_5 U$$4292/B input215/X dadda_fa_1_62_5/CIN VGND VGND VPWR VPWR dadda_fa_2_63_2/A
+ dadda_fa_2_62_5/A sky130_fd_sc_hd__fa_1
XFILLER_87_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_55_4 U$$2378/X U$$2511/X U$$2644/X VGND VGND VPWR VPWR dadda_fa_2_56_1/CIN
+ dadda_fa_2_55_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_48_3 U$$1300/X U$$1433/X U$$1566/X VGND VGND VPWR VPWR dadda_fa_2_49_2/A
+ dadda_fa_2_48_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_25_2 dadda_fa_4_25_2/A dadda_fa_4_25_2/B dadda_fa_4_25_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_26_0/CIN dadda_fa_5_25_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_18_1 input166/X dadda_fa_4_18_1/B dadda_fa_4_18_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_5_19_0/B dadda_fa_5_18_1/B sky130_fd_sc_hd__fa_1
XFILLER_169_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1603 U$$2862/B1 VGND VGND VPWR VPWR U$$2042/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1614 U$$4506/A1 VGND VGND VPWR VPWR U$$4367/B1 sky130_fd_sc_hd__buf_4
XFILLER_104_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1625 U$$4504/A1 VGND VGND VPWR VPWR U$$4093/A1 sky130_fd_sc_hd__buf_2
Xfanout1636 input115/X VGND VGND VPWR VPWR U$$2993/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1647 U$$2578/B1 VGND VGND VPWR VPWR U$$388/A1 sky130_fd_sc_hd__buf_6
Xfanout660 U$$902/B2 VGND VGND VPWR VPWR U$$898/B2 sky130_fd_sc_hd__buf_4
XU$$4106 U$$4106/A U$$4108/B VGND VGND VPWR VPWR U$$4106/X sky130_fd_sc_hd__xor2_1
Xfanout1658 U$$2578/A1 VGND VGND VPWR VPWR U$$384/B1 sky130_fd_sc_hd__buf_2
Xfanout671 U$$690/X VGND VGND VPWR VPWR U$$807/B2 sky130_fd_sc_hd__buf_4
Xdadda_ha_3_21_3 U$$1246/X U$$1379/X VGND VGND VPWR VPWR dadda_fa_4_22_1/B dadda_ha_3_21_3/SUM
+ sky130_fd_sc_hd__ha_1
Xfanout1669 U$$4494/A1 VGND VGND VPWR VPWR U$$4081/B1 sky130_fd_sc_hd__buf_4
XU$$4117 U$$4117/A U$$4133/B VGND VGND VPWR VPWR U$$4117/X sky130_fd_sc_hd__xor2_1
XFILLER_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4128 U$$4400/B1 U$$4158/A2 U$$4265/B1 U$$4158/B2 VGND VGND VPWR VPWR U$$4129/A
+ sky130_fd_sc_hd__a22o_1
Xfanout682 U$$642/B2 VGND VGND VPWR VPWR U$$682/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout693 U$$543/B2 VGND VGND VPWR VPWR U$$497/B2 sky130_fd_sc_hd__buf_4
XU$$4139 U$$4139/A U$$4159/B VGND VGND VPWR VPWR U$$4139/X sky130_fd_sc_hd__xor2_1
XU$$3405 U$$3405/A U$$3411/B VGND VGND VPWR VPWR U$$3405/X sky130_fd_sc_hd__xor2_1
XFILLER_19_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3416 U$$3416/A1 U$$3416/A2 U$$3418/A1 U$$3416/B2 VGND VGND VPWR VPWR U$$3417/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3427 U$$3562/A VGND VGND VPWR VPWR U$$3427/Y sky130_fd_sc_hd__inv_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3438 U$$3438/A U$$3482/B VGND VGND VPWR VPWR U$$3438/X sky130_fd_sc_hd__xor2_1
XU$$2704 U$$2704/A U$$2708/B VGND VGND VPWR VPWR U$$2704/X sky130_fd_sc_hd__xor2_1
XU$$3449 U$$4132/B1 U$$3473/A2 U$$3999/A1 U$$3473/B2 VGND VGND VPWR VPWR U$$3450/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2715 U$$4220/B1 U$$2733/A2 U$$4361/A1 U$$2733/B2 VGND VGND VPWR VPWR U$$2716/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2726 U$$2726/A U$$2738/B VGND VGND VPWR VPWR U$$2726/X sky130_fd_sc_hd__xor2_1
XU$$2737 U$$3285/A1 U$$2737/A2 U$$2737/B1 U$$2737/B2 VGND VGND VPWR VPWR U$$2738/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2748 U$$2748/A1 U$$2804/A2 U$$4257/A1 U$$2804/B2 VGND VGND VPWR VPWR U$$2749/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_1 U$$446/X U$$579/X U$$712/X VGND VGND VPWR VPWR dadda_fa_4_21_0/CIN
+ dadda_fa_4_20_2/A sky130_fd_sc_hd__fa_1
XU$$2759 U$$2759/A U$$2799/B VGND VGND VPWR VPWR U$$2759/X sky130_fd_sc_hd__xor2_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_416_ _416_/CLK _416_/D VGND VGND VPWR VPWR _416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_347_ _349_/CLK _347_/D VGND VGND VPWR VPWR _347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_278_ _408_/CLK _278_/D VGND VGND VPWR VPWR _278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_100_0_1931 VGND VGND VPWR VPWR dadda_fa_2_100_0/A dadda_fa_2_100_0_1931/LO
+ sky130_fd_sc_hd__conb_1
Xdadda_fa_2_72_4 dadda_fa_2_72_4/A dadda_fa_2_72_4/B dadda_fa_2_72_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_1/CIN dadda_fa_3_72_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_65_3 dadda_fa_2_65_3/A dadda_fa_2_65_3/B dadda_fa_2_65_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_1/B dadda_fa_3_65_3/B sky130_fd_sc_hd__fa_1
XFILLER_110_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_58_2 dadda_fa_2_58_2/A dadda_fa_2_58_2/B dadda_fa_2_58_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_1/A dadda_fa_3_58_3/A sky130_fd_sc_hd__fa_1
XFILLER_77_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_35_1 dadda_fa_5_35_1/A dadda_fa_5_35_1/B dadda_fa_5_35_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_36_0/B dadda_fa_7_35_0/A sky130_fd_sc_hd__fa_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_28_0 dadda_fa_5_28_0/A dadda_fa_5_28_0/B dadda_fa_5_28_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_29_0/A dadda_fa_6_28_0/CIN sky130_fd_sc_hd__fa_1
XU$$3950 U$$4361/A1 U$$3970/A2 U$$4363/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3951/A
+ sky130_fd_sc_hd__a22o_1
XU$$3961 U$$3961/A U$$3961/B VGND VGND VPWR VPWR U$$3961/X sky130_fd_sc_hd__xor2_1
XFILLER_65_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3972 U$$3972/A VGND VGND VPWR VPWR U$$3972/Y sky130_fd_sc_hd__inv_1
XU$$3983 U$$4257/A1 U$$4025/A2 U$$4257/B1 U$$4025/B2 VGND VGND VPWR VPWR U$$3984/A
+ sky130_fd_sc_hd__a22o_1
XU$$3994 U$$3994/A U$$4026/B VGND VGND VPWR VPWR U$$3994/X sky130_fd_sc_hd__xor2_1
XFILLER_91_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_88_0_1927 VGND VGND VPWR VPWR dadda_fa_1_88_0/A dadda_fa_1_88_0_1927/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_118_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_102_0 dadda_fa_5_102_0/A dadda_fa_5_102_0/B dadda_fa_5_102_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_103_0/A dadda_fa_6_102_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_145_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput263 output263/A VGND VGND VPWR VPWR o[105] sky130_fd_sc_hd__buf_2
Xoutput274 output274/A VGND VGND VPWR VPWR o[115] sky130_fd_sc_hd__buf_2
XFILLER_87_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput285 output285/A VGND VGND VPWR VPWR o[125] sky130_fd_sc_hd__buf_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput296 output296/A VGND VGND VPWR VPWR o[1] sky130_fd_sc_hd__buf_2
XFILLER_87_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_60_2 U$$2787/X U$$2920/X U$$3053/X VGND VGND VPWR VPWR dadda_fa_2_61_1/A
+ dadda_fa_2_60_4/A sky130_fd_sc_hd__fa_1
XFILLER_47_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_831 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_1 U$$778/X U$$911/X U$$1044/X VGND VGND VPWR VPWR dadda_fa_2_54_0/CIN
+ dadda_fa_2_53_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_4_30_0 dadda_fa_4_30_0/A dadda_fa_4_30_0/B dadda_fa_4_30_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_31_0/A dadda_fa_5_30_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_46_0 U$$99/X U$$232/X U$$365/X VGND VGND VPWR VPWR dadda_fa_2_47_1/CIN
+ dadda_fa_2_46_4/A sky130_fd_sc_hd__fa_1
XFILLER_82_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_201_ _201_/CLK _201_/D VGND VGND VPWR VPWR _201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1104 final_adder.U$$174/A final_adder.U$$883/X VGND VGND VPWR VPWR
+ output363/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1115 final_adder.U$$164/B final_adder.U$$935/X VGND VGND VPWR VPWR
+ output375/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1126 final_adder.U$$152/A final_adder.U$$861/X VGND VGND VPWR VPWR
+ output260/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1137 final_adder.U$$142/B final_adder.U$$913/X VGND VGND VPWR VPWR
+ output272/A sky130_fd_sc_hd__xor2_1
XFILLER_137_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1148 final_adder.U$$130/A final_adder.U$$839/X VGND VGND VPWR VPWR
+ output284/A sky130_fd_sc_hd__xor2_1
XFILLER_171_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_82_3 dadda_fa_3_82_3/A dadda_fa_3_82_3/B dadda_fa_3_82_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_1/B dadda_fa_4_82_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_75_2 dadda_fa_3_75_2/A dadda_fa_3_75_2/B dadda_fa_3_75_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_1/A dadda_fa_4_75_2/B sky130_fd_sc_hd__fa_1
XFILLER_78_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1400 U$$254/B VGND VGND VPWR VPWR U$$210/B sky130_fd_sc_hd__buf_4
Xfanout1411 U$$2541/B VGND VGND VPWR VPWR U$$2529/B sky130_fd_sc_hd__buf_6
Xdadda_fa_3_68_1 dadda_fa_3_68_1/A dadda_fa_3_68_1/B dadda_fa_3_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_0/CIN dadda_fa_4_68_2/A sky130_fd_sc_hd__fa_1
Xfanout1422 U$$822/A VGND VGND VPWR VPWR U$$804/B sky130_fd_sc_hd__buf_4
XFILLER_120_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_45_0 dadda_fa_6_45_0/A dadda_fa_6_45_0/B dadda_fa_6_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_46_0/B dadda_fa_7_45_0/CIN sky130_fd_sc_hd__fa_1
Xfanout1433 fanout1438/X VGND VGND VPWR VPWR U$$2408/B sky130_fd_sc_hd__buf_4
Xfanout1444 U$$2301/B VGND VGND VPWR VPWR U$$2329/A sky130_fd_sc_hd__clkbuf_8
Xfanout1455 U$$2186/B VGND VGND VPWR VPWR U$$2168/B sky130_fd_sc_hd__buf_6
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1466 U$$2054/A VGND VGND VPWR VPWR U$$2053/B sky130_fd_sc_hd__buf_8
Xfanout1477 U$$1727/B VGND VGND VPWR VPWR U$$1697/B sky130_fd_sc_hd__buf_6
XFILLER_66_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout490 U$$3557/A2 VGND VGND VPWR VPWR U$$3559/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout1488 U$$1618/B VGND VGND VPWR VPWR U$$1594/B sky130_fd_sc_hd__clkbuf_4
XU$$3202 U$$3202/A U$$3208/B VGND VGND VPWR VPWR U$$3202/X sky130_fd_sc_hd__xor2_1
Xfanout1499 U$$1449/B VGND VGND VPWR VPWR U$$1415/B sky130_fd_sc_hd__buf_6
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3213 U$$4446/A1 U$$3255/A2 U$$4446/B1 U$$3255/B2 VGND VGND VPWR VPWR U$$3214/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3224 U$$3224/A U$$3242/B VGND VGND VPWR VPWR U$$3224/X sky130_fd_sc_hd__xor2_1
XU$$3235 U$$3370/B1 U$$3241/A2 U$$3372/B1 U$$3241/B2 VGND VGND VPWR VPWR U$$3236/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$17 _313_/Q _185_/Q VGND VGND VPWR VPWR final_adder.U$$239/B1 final_adder.U$$238/B
+ sky130_fd_sc_hd__ha_1
XFILLER_62_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2501 U$$2501/A U$$2545/B VGND VGND VPWR VPWR U$$2501/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$28 _324_/Q _196_/Q VGND VGND VPWR VPWR final_adder.U$$997/B1 final_adder.U$$226/A
+ sky130_fd_sc_hd__ha_1
XU$$3246 U$$3246/A U$$3288/A VGND VGND VPWR VPWR U$$3246/X sky130_fd_sc_hd__xor2_1
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2512 U$$46/A1 U$$2546/A2 U$$48/A1 U$$2546/B2 VGND VGND VPWR VPWR U$$2513/A sky130_fd_sc_hd__a22o_1
XU$$3257 U$$517/A1 U$$3257/A2 U$$517/B1 U$$3257/B2 VGND VGND VPWR VPWR U$$3258/A sky130_fd_sc_hd__a22o_1
XU$$3268 U$$3268/A U$$3284/B VGND VGND VPWR VPWR U$$3268/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$39 _335_/Q _207_/Q VGND VGND VPWR VPWR final_adder.U$$217/B1 final_adder.U$$216/B
+ sky130_fd_sc_hd__ha_1
XU$$2523 U$$2523/A U$$2529/B VGND VGND VPWR VPWR U$$2523/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_104_2 dadda_fa_4_104_2/A dadda_fa_4_104_2/B dadda_fa_4_104_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_105_0/CIN dadda_fa_5_104_1/CIN sky130_fd_sc_hd__fa_1
XU$$2534 U$$3628/B1 U$$2540/A2 U$$3630/B1 U$$2540/B2 VGND VGND VPWR VPWR U$$2535/A
+ sky130_fd_sc_hd__a22o_1
XU$$3279 U$$3416/A1 U$$3283/A2 U$$3418/A1 U$$3283/B2 VGND VGND VPWR VPWR U$$3280/A
+ sky130_fd_sc_hd__a22o_1
XU$$1800 U$$1800/A U$$1836/B VGND VGND VPWR VPWR U$$1800/X sky130_fd_sc_hd__xor2_1
XU$$2545 U$$2545/A U$$2545/B VGND VGND VPWR VPWR U$$2545/X sky130_fd_sc_hd__xor2_1
XFILLER_62_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$2556 U$$3650/B1 U$$2574/A2 U$$3515/B1 U$$2574/B2 VGND VGND VPWR VPWR U$$2557/A
+ sky130_fd_sc_hd__a22o_1
XU$$1811 U$$576/B1 U$$1841/A2 U$$443/A1 U$$1841/B2 VGND VGND VPWR VPWR U$$1812/A sky130_fd_sc_hd__a22o_1
XU$$1822 U$$1822/A U$$1828/B VGND VGND VPWR VPWR U$$1822/X sky130_fd_sc_hd__xor2_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2567 U$$2567/A U$$2575/B VGND VGND VPWR VPWR U$$2567/X sky130_fd_sc_hd__xor2_1
XFILLER_61_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1833 U$$52/A1 U$$1841/A2 U$$54/A1 U$$1841/B2 VGND VGND VPWR VPWR U$$1834/A sky130_fd_sc_hd__a22o_1
XU$$2578 U$$2578/A1 U$$2578/A2 U$$2578/B1 U$$2578/B2 VGND VGND VPWR VPWR U$$2579/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2589 U$$2589/A U$$2591/B VGND VGND VPWR VPWR U$$2589/X sky130_fd_sc_hd__xor2_1
XU$$1844 U$$1844/A U$$1854/B VGND VGND VPWR VPWR U$$1844/X sky130_fd_sc_hd__xor2_1
XU$$1855 U$$620/B1 U$$1859/A2 U$$898/A1 U$$1859/B2 VGND VGND VPWR VPWR U$$1856/A sky130_fd_sc_hd__a22o_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1866 U$$1866/A U$$1874/B VGND VGND VPWR VPWR U$$1866/X sky130_fd_sc_hd__xor2_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1877 U$$918/A1 U$$1915/A2 U$$920/A1 U$$1915/B2 VGND VGND VPWR VPWR U$$1878/A sky130_fd_sc_hd__a22o_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1888 U$$1888/A U$$1916/B VGND VGND VPWR VPWR U$$1888/X sky130_fd_sc_hd__xor2_1
XFILLER_148_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1899 U$$2310/A1 U$$1911/A2 U$$942/A1 U$$1911/B2 VGND VGND VPWR VPWR U$$1900/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_118_0 dadda_fa_7_118_0/A dadda_fa_7_118_0/B dadda_fa_7_118_0/CIN VGND
+ VGND VPWR VPWR _415_/D _286_/D sky130_fd_sc_hd__fa_1
XFILLER_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_76_0_1922 VGND VGND VPWR VPWR dadda_fa_0_76_0/A dadda_fa_0_76_0_1922/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_147_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_70_1 dadda_fa_2_70_1/A dadda_fa_2_70_1/B dadda_fa_2_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_0/CIN dadda_fa_3_70_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_63_0 dadda_fa_2_63_0/A dadda_fa_2_63_0/B dadda_fa_2_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_0/B dadda_fa_3_63_2/B sky130_fd_sc_hd__fa_1
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$518 final_adder.U$$526/B final_adder.U$$518/B VGND VGND VPWR VPWR
+ final_adder.U$$638/B sky130_fd_sc_hd__and2_1
XFILLER_97_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$529 final_adder.U$$528/B final_adder.U$$413/X final_adder.U$$405/X
+ VGND VGND VPWR VPWR final_adder.U$$529/X sky130_fd_sc_hd__a21o_1
XFILLER_111_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$4470 U$$4470/A1 U$$4388/X U$$4472/A1 U$$4492/B2 VGND VGND VPWR VPWR U$$4471/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4481 U$$4481/A U$$4481/B VGND VGND VPWR VPWR U$$4481/X sky130_fd_sc_hd__xor2_1
XU$$4492 U$$4492/A1 U$$4388/X U$$4492/B1 U$$4492/B2 VGND VGND VPWR VPWR U$$4493/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$3780 U$$3780/A U$$3828/B VGND VGND VPWR VPWR U$$3780/X sky130_fd_sc_hd__xor2_1
XU$$3791 U$$4476/A1 U$$3791/A2 U$$4478/A1 U$$3791/B2 VGND VGND VPWR VPWR U$$3792/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_92_2 dadda_fa_4_92_2/A dadda_fa_4_92_2/B dadda_fa_4_92_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_93_0/CIN dadda_fa_5_92_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_4_85_1 dadda_fa_4_85_1/A dadda_fa_4_85_1/B dadda_fa_4_85_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_86_0/B dadda_fa_5_85_1/B sky130_fd_sc_hd__fa_1
XFILLER_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_7_62_0 dadda_fa_7_62_0/A dadda_fa_7_62_0/B dadda_fa_7_62_0/CIN VGND VGND
+ VPWR VPWR _359_/D _230_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_78_0 dadda_fa_4_78_0/A dadda_fa_4_78_0/B dadda_fa_4_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_79_0/A dadda_fa_5_78_1/A sky130_fd_sc_hd__fa_1
XFILLER_134_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$902 U$$902/A1 U$$902/A2 U$$902/B1 U$$902/B2 VGND VGND VPWR VPWR U$$903/A sky130_fd_sc_hd__a22o_1
XFILLER_91_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$913 U$$913/A U$$913/B VGND VGND VPWR VPWR U$$913/X sky130_fd_sc_hd__xor2_1
XU$$924 U$$924/A1 U$$942/A2 U$$926/A1 U$$942/B2 VGND VGND VPWR VPWR U$$925/A sky130_fd_sc_hd__a22o_1
XFILLER_84_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$935 U$$935/A U$$959/A VGND VGND VPWR VPWR U$$935/X sky130_fd_sc_hd__xor2_1
XU$$946 U$$946/A1 U$$956/A2 U$$948/A1 U$$956/B2 VGND VGND VPWR VPWR U$$947/A sky130_fd_sc_hd__a22o_1
XFILLER_56_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$957 U$$957/A U$$958/A VGND VGND VPWR VPWR U$$957/X sky130_fd_sc_hd__xor2_1
XU$$968 U$$968/A U$$982/B VGND VGND VPWR VPWR U$$968/X sky130_fd_sc_hd__xor2_1
XU$$1107 U$$1107/A U$$1175/B VGND VGND VPWR VPWR U$$1107/X sky130_fd_sc_hd__xor2_1
XFILLER_141_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1118 U$$2897/B1 U$$1194/A2 U$$981/B1 U$$1194/B2 VGND VGND VPWR VPWR U$$1119/A
+ sky130_fd_sc_hd__a22o_1
XU$$979 U$$979/A1 U$$979/A2 U$$979/B1 U$$979/B2 VGND VGND VPWR VPWR U$$980/A sky130_fd_sc_hd__a22o_1
XU$$1129 U$$1129/A U$$1163/B VGND VGND VPWR VPWR U$$1129/X sky130_fd_sc_hd__xor2_1
XFILLER_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_80_0 dadda_fa_3_80_0/A dadda_fa_3_80_0/B dadda_fa_3_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_0/B dadda_fa_4_80_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_112_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1230 U$$3314/B1 VGND VGND VPWR VPWR U$$576/A1 sky130_fd_sc_hd__buf_4
XFILLER_67_926 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1241 U$$3979/B1 VGND VGND VPWR VPWR U$$967/A1 sky130_fd_sc_hd__buf_4
XFILLER_121_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1252 U$$547/A VGND VGND VPWR VPWR U$$498/B sky130_fd_sc_hd__buf_6
Xfanout1263 input60/X VGND VGND VPWR VPWR U$$4384/A sky130_fd_sc_hd__buf_6
Xfanout1274 U$$4191/B VGND VGND VPWR VPWR U$$4231/B sky130_fd_sc_hd__buf_6
Xfanout1285 U$$341/B VGND VGND VPWR VPWR U$$313/B sky130_fd_sc_hd__buf_4
Xfanout1296 U$$4058/B VGND VGND VPWR VPWR U$$4082/B sky130_fd_sc_hd__buf_6
XU$$3010 U$$3010/A U$$3013/A VGND VGND VPWR VPWR U$$3010/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_42_5 dadda_fa_2_42_5/A dadda_fa_2_42_5/B dadda_fa_2_42_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_43_2/A dadda_fa_4_42_0/A sky130_fd_sc_hd__fa_2
XU$$3021 U$$3021/A U$$3061/B VGND VGND VPWR VPWR U$$3021/X sky130_fd_sc_hd__xor2_1
XFILLER_75_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3032 U$$840/A1 U$$3124/A2 U$$840/B1 U$$3124/B2 VGND VGND VPWR VPWR U$$3033/A sky130_fd_sc_hd__a22o_1
XFILLER_75_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3043 U$$3043/A U$$3077/B VGND VGND VPWR VPWR U$$3043/X sky130_fd_sc_hd__xor2_1
XU$$3054 U$$3189/B1 U$$3066/A2 U$$3056/A1 U$$3066/B2 VGND VGND VPWR VPWR U$$3055/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3065 U$$3065/A U$$3073/B VGND VGND VPWR VPWR U$$3065/X sky130_fd_sc_hd__xor2_1
XU$$2320 U$$3964/A1 U$$2320/A2 U$$3966/A1 U$$2320/B2 VGND VGND VPWR VPWR U$$2321/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_35_4 U$$1939/X U$$2072/X U$$2205/X VGND VGND VPWR VPWR dadda_fa_3_36_1/CIN
+ dadda_fa_3_35_3/CIN sky130_fd_sc_hd__fa_1
XU$$2331 U$$2446/B VGND VGND VPWR VPWR U$$2331/Y sky130_fd_sc_hd__inv_1
XU$$3076 U$$745/B1 U$$3124/A2 U$$612/A1 U$$3124/B2 VGND VGND VPWR VPWR U$$3077/A sky130_fd_sc_hd__a22o_1
XU$$2342 U$$2342/A U$$2412/B VGND VGND VPWR VPWR U$$2342/X sky130_fd_sc_hd__xor2_1
XU$$3087 U$$3087/A U$$3119/B VGND VGND VPWR VPWR U$$3087/X sky130_fd_sc_hd__xor2_1
XU$$2353 U$$983/A1 U$$2395/A2 U$$983/B1 U$$2395/B2 VGND VGND VPWR VPWR U$$2354/A sky130_fd_sc_hd__a22o_1
XU$$3098 U$$3370/B1 U$$3108/A2 U$$3372/B1 U$$3108/B2 VGND VGND VPWR VPWR U$$3099/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2364 U$$2364/A U$$2402/B VGND VGND VPWR VPWR U$$2364/X sky130_fd_sc_hd__xor2_1
XU$$1630 U$$1630/A U$$1630/B VGND VGND VPWR VPWR U$$1630/X sky130_fd_sc_hd__xor2_1
XU$$2375 U$$183/A1 U$$2413/A2 U$$870/A1 U$$2413/B2 VGND VGND VPWR VPWR U$$2376/A sky130_fd_sc_hd__a22o_1
XU$$1641 U$$4244/A1 U$$1641/A2 U$$1641/B1 U$$1641/B2 VGND VGND VPWR VPWR U$$1642/A
+ sky130_fd_sc_hd__a22o_1
XU$$2386 U$$2386/A U$$2402/B VGND VGND VPWR VPWR U$$2386/X sky130_fd_sc_hd__xor2_1
XU$$2397 U$$3628/B1 U$$2407/A2 U$$70/A1 U$$2407/B2 VGND VGND VPWR VPWR U$$2398/A sky130_fd_sc_hd__a22o_1
XU$$1652 U$$2748/A1 U$$1698/A2 U$$3296/B1 U$$1698/B2 VGND VGND VPWR VPWR U$$1653/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1663 U$$1663/A U$$1699/B VGND VGND VPWR VPWR U$$1663/X sky130_fd_sc_hd__xor2_1
XU$$1674 U$$30/A1 U$$1702/A2 U$$32/A1 U$$1702/B2 VGND VGND VPWR VPWR U$$1675/A sky130_fd_sc_hd__a22o_1
XU$$1685 U$$1685/A U$$1699/B VGND VGND VPWR VPWR U$$1685/X sky130_fd_sc_hd__xor2_1
XU$$1696 U$$52/A1 U$$1696/A2 U$$54/A1 U$$1696/B2 VGND VGND VPWR VPWR U$$1697/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_95_0 dadda_fa_5_95_0/A dadda_fa_5_95_0/B dadda_fa_5_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_96_0/A dadda_fa_6_95_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$304 final_adder.U$$306/B final_adder.U$$304/B VGND VGND VPWR VPWR
+ final_adder.U$$430/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$315 final_adder.U$$314/B final_adder.U$$189/X final_adder.U$$187/X
+ VGND VGND VPWR VPWR final_adder.U$$315/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$326 final_adder.U$$328/B final_adder.U$$326/B VGND VGND VPWR VPWR
+ final_adder.U$$452/B sky130_fd_sc_hd__and2_1
XFILLER_111_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$337 final_adder.U$$336/B final_adder.U$$211/X final_adder.U$$209/X
+ VGND VGND VPWR VPWR final_adder.U$$337/X sky130_fd_sc_hd__a21o_1
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$348 final_adder.U$$350/B final_adder.U$$348/B VGND VGND VPWR VPWR
+ final_adder.U$$474/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$359 final_adder.U$$358/B final_adder.U$$233/X final_adder.U$$231/X
+ VGND VGND VPWR VPWR final_adder.U$$359/X sky130_fd_sc_hd__a21o_1
XU$$209 U$$72/A1 U$$213/A2 U$$74/A1 U$$213/B2 VGND VGND VPWR VPWR U$$210/A sky130_fd_sc_hd__a22o_1
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_111_2 U$$4086/X U$$4219/X U$$4352/X VGND VGND VPWR VPWR dadda_fa_4_112_1/CIN
+ dadda_fa_4_111_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_104_1 U$$4205/X U$$4338/X U$$4471/X VGND VGND VPWR VPWR dadda_fa_4_105_0/CIN
+ dadda_fa_4_104_2/A sky130_fd_sc_hd__fa_1
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_6_125_0 input157/X dadda_fa_6_125_0/B dadda_fa_6_125_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_126_0/B dadda_fa_7_125_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_68_4 U$$1872/X U$$2005/X U$$2138/X VGND VGND VPWR VPWR dadda_fa_1_69_7/A
+ dadda_fa_1_68_8/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_45_3 dadda_fa_3_45_3/A dadda_fa_3_45_3/B dadda_fa_3_45_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_1/B dadda_fa_4_45_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$871 final_adder.U$$774/X final_adder.U$$727/X final_adder.U$$775/X
+ VGND VGND VPWR VPWR final_adder.U$$871/X sky130_fd_sc_hd__a21o_1
XFILLER_91_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$710 U$$710/A U$$744/B VGND VGND VPWR VPWR U$$710/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_38_2 dadda_fa_3_38_2/A dadda_fa_3_38_2/B dadda_fa_3_38_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_1/A dadda_fa_4_38_2/B sky130_fd_sc_hd__fa_1
XFILLER_16_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$721 U$$721/A1 U$$769/A2 U$$721/B1 U$$769/B2 VGND VGND VPWR VPWR U$$722/A sky130_fd_sc_hd__a22o_1
XFILLER_63_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$893 final_adder.U$$796/X final_adder.U$$505/X final_adder.U$$797/X
+ VGND VGND VPWR VPWR final_adder.U$$893/X sky130_fd_sc_hd__a21o_1
XU$$732 U$$732/A U$$768/B VGND VGND VPWR VPWR U$$732/X sky130_fd_sc_hd__xor2_1
XU$$743 U$$878/B1 U$$743/A2 U$$745/A1 U$$743/B2 VGND VGND VPWR VPWR U$$744/A sky130_fd_sc_hd__a22o_1
XFILLER_16_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$754 U$$754/A U$$768/B VGND VGND VPWR VPWR U$$754/X sky130_fd_sc_hd__xor2_1
XU$$765 U$$900/B1 U$$809/A2 U$$765/B1 U$$809/B2 VGND VGND VPWR VPWR U$$766/A sky130_fd_sc_hd__a22o_1
XFILLER_90_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$776 U$$776/A U$$778/B VGND VGND VPWR VPWR U$$776/X sky130_fd_sc_hd__xor2_1
XFILLER_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$787 U$$787/A1 U$$817/A2 U$$787/B1 U$$817/B2 VGND VGND VPWR VPWR U$$788/A sky130_fd_sc_hd__a22o_1
XFILLER_16_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XU$$798 U$$798/A U$$804/B VGND VGND VPWR VPWR U$$798/X sky130_fd_sc_hd__xor2_1
XFILLER_71_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1060 U$$3080/A1 VGND VGND VPWR VPWR U$$4450/A1 sky130_fd_sc_hd__clkbuf_8
Xdadda_ha_2_27_2 U$$859/X U$$992/X VGND VGND VPWR VPWR dadda_fa_3_28_2/CIN dadda_fa_4_27_0/A
+ sky130_fd_sc_hd__ha_1
Xfanout1071 U$$2665/A1 VGND VGND VPWR VPWR U$$884/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1082 input83/X VGND VGND VPWR VPWR U$$745/A1 sky130_fd_sc_hd__buf_6
Xfanout1093 input82/X VGND VGND VPWR VPWR U$$3618/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_54_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_40_2 U$$2348/X U$$2481/X U$$2614/X VGND VGND VPWR VPWR dadda_fa_3_41_1/A
+ dadda_fa_3_40_3/A sky130_fd_sc_hd__fa_1
XFILLER_82_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_33_1 U$$472/X U$$605/X U$$738/X VGND VGND VPWR VPWR dadda_fa_3_34_0/CIN
+ dadda_fa_3_33_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2150 U$$2150/A U$$2191/A VGND VGND VPWR VPWR U$$2150/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_10_0 U$$692/X U$$778/B input140/X VGND VGND VPWR VPWR dadda_fa_6_11_0/A
+ dadda_fa_6_10_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_26_0 U$$59/X U$$192/X U$$325/X VGND VGND VPWR VPWR dadda_fa_3_27_2/B dadda_fa_3_26_3/B
+ sky130_fd_sc_hd__fa_1
XU$$2161 U$$2844/B1 U$$2177/A2 U$$2574/A1 U$$2177/B2 VGND VGND VPWR VPWR U$$2162/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2172 U$$2172/A U$$2192/A VGND VGND VPWR VPWR U$$2172/X sky130_fd_sc_hd__xor2_1
XU$$2183 U$$2183/A1 U$$2189/A2 U$$4512/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2184/A
+ sky130_fd_sc_hd__a22o_1
XU$$2194 U$$2329/A VGND VGND VPWR VPWR U$$2194/Y sky130_fd_sc_hd__inv_1
XU$$1460 U$$90/A1 U$$1460/A2 U$$92/A1 U$$1460/B2 VGND VGND VPWR VPWR U$$1461/A sky130_fd_sc_hd__a22o_1
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1471 U$$1471/A U$$1497/B VGND VGND VPWR VPWR U$$1471/X sky130_fd_sc_hd__xor2_1
XU$$1482 U$$521/B1 U$$1502/A2 U$$386/B1 U$$1502/B2 VGND VGND VPWR VPWR U$$1483/A sky130_fd_sc_hd__a22o_1
XU$$1493 U$$1493/A input14/X VGND VGND VPWR VPWR U$$1493/X sky130_fd_sc_hd__xor2_1
XFILLER_124_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_85_4 U$$3103/X U$$3236/X U$$3369/X VGND VGND VPWR VPWR dadda_fa_2_86_3/CIN
+ dadda_fa_2_85_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_131_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_78_3 U$$2424/X U$$2557/X U$$2690/X VGND VGND VPWR VPWR dadda_fa_2_79_1/B
+ dadda_fa_2_78_4/B sky130_fd_sc_hd__fa_1
XFILLER_44_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_55_2 dadda_fa_4_55_2/A dadda_fa_4_55_2/B dadda_fa_4_55_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_56_0/CIN dadda_fa_5_55_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$101 _397_/Q _269_/Q VGND VGND VPWR VPWR final_adder.U$$155/B1 final_adder.U$$154/B
+ sky130_fd_sc_hd__ha_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$112 _408_/Q _280_/Q VGND VGND VPWR VPWR final_adder.U$$913/B1 final_adder.U$$142/A
+ sky130_fd_sc_hd__ha_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_48_1 dadda_fa_4_48_1/A dadda_fa_4_48_1/B dadda_fa_4_48_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_49_0/B dadda_fa_5_48_1/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$123 _419_/Q _291_/Q VGND VGND VPWR VPWR final_adder.U$$133/B1 final_adder.U$$132/B
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$134 final_adder.U$$134/A final_adder.U$$134/B VGND VGND VPWR VPWR
+ final_adder.U$$262/B sky130_fd_sc_hd__and2_1
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$145 final_adder.U$$144/B final_adder.U$$915/B1 final_adder.U$$145/B1
+ VGND VGND VPWR VPWR final_adder.U$$145/X sky130_fd_sc_hd__a21o_1
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_25_0 dadda_fa_7_25_0/A dadda_fa_7_25_0/B dadda_fa_7_25_0/CIN VGND VGND
+ VPWR VPWR _322_/D _193_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$156 final_adder.U$$156/A final_adder.U$$156/B VGND VGND VPWR VPWR
+ final_adder.U$$284/B sky130_fd_sc_hd__and2_1
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$167 final_adder.U$$166/B final_adder.U$$937/B1 final_adder.U$$167/B1
+ VGND VGND VPWR VPWR final_adder.U$$167/X sky130_fd_sc_hd__a21o_2
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$178 final_adder.U$$178/A final_adder.U$$178/B VGND VGND VPWR VPWR
+ final_adder.U$$306/B sky130_fd_sc_hd__and2_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$189 final_adder.U$$188/B final_adder.U$$959/B1 final_adder.U$$189/B1
+ VGND VGND VPWR VPWR final_adder.U$$189/X sky130_fd_sc_hd__a21o_1
XFILLER_57_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_380_ _380_/CLK _380_/D VGND VGND VPWR VPWR _380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_0_73_2 U$$1483/X U$$1616/X U$$1749/X VGND VGND VPWR VPWR dadda_fa_1_74_8/A
+ dadda_fa_2_73_0/A sky130_fd_sc_hd__fa_1
XFILLER_95_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput130 c[100] VGND VGND VPWR VPWR input130/X sky130_fd_sc_hd__clkbuf_4
XFILLER_163_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput141 c[110] VGND VGND VPWR VPWR input141/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_3_50_1 dadda_fa_3_50_1/A dadda_fa_3_50_1/B dadda_fa_3_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_0/CIN dadda_fa_4_50_2/A sky130_fd_sc_hd__fa_1
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_66_1 U$$538/X U$$671/X U$$804/X VGND VGND VPWR VPWR dadda_fa_1_67_5/CIN
+ dadda_fa_1_66_7/CIN sky130_fd_sc_hd__fa_1
Xinput152 c[120] VGND VGND VPWR VPWR input152/X sky130_fd_sc_hd__buf_2
Xinput163 c[15] VGND VGND VPWR VPWR input163/X sky130_fd_sc_hd__buf_2
XFILLER_76_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_3_43_0 dadda_fa_3_43_0/A dadda_fa_3_43_0/B dadda_fa_3_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_0/B dadda_fa_4_43_1/CIN sky130_fd_sc_hd__fa_1
Xinput174 c[25] VGND VGND VPWR VPWR input174/X sky130_fd_sc_hd__clkbuf_2
Xinput185 c[35] VGND VGND VPWR VPWR input185/X sky130_fd_sc_hd__clkbuf_4
XFILLER_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput196 c[45] VGND VGND VPWR VPWR input196/X sky130_fd_sc_hd__dlymetal6s2s_1
Xdadda_fa_0_59_0 U$$125/X U$$258/X U$$391/X VGND VGND VPWR VPWR dadda_fa_1_60_6/B
+ dadda_fa_1_59_8/A sky130_fd_sc_hd__fa_2
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$690 final_adder.U$$706/B final_adder.U$$690/B VGND VGND VPWR VPWR
+ final_adder.U$$770/A sky130_fd_sc_hd__and2_1
XFILLER_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$540 U$$540/A U$$548/A VGND VGND VPWR VPWR U$$540/X sky130_fd_sc_hd__xor2_1
XFILLER_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$551 U$$669/B U$$551/B VGND VGND VPWR VPWR U$$551/X sky130_fd_sc_hd__and2_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$562 U$$562/A1 U$$642/A2 U$$562/B1 U$$642/B2 VGND VGND VPWR VPWR U$$563/A sky130_fd_sc_hd__a22o_1
XU$$573 U$$573/A U$$639/B VGND VGND VPWR VPWR U$$573/X sky130_fd_sc_hd__xor2_1
XU$$584 U$$721/A1 U$$636/A2 U$$721/B1 U$$636/B2 VGND VGND VPWR VPWR U$$585/A sky130_fd_sc_hd__a22o_1
XFILLER_72_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$595 U$$595/A U$$631/B VGND VGND VPWR VPWR U$$595/X sky130_fd_sc_hd__xor2_1
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_100_0 dadda_fa_7_100_0/A dadda_fa_7_100_0/B dadda_fa_7_100_0/CIN VGND
+ VGND VPWR VPWR _397_/D _268_/D sky130_fd_sc_hd__fa_1
XFILLER_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_95_3 U$$3788/X U$$3921/X U$$4054/X VGND VGND VPWR VPWR dadda_fa_3_96_1/B
+ dadda_fa_3_95_3/B sky130_fd_sc_hd__fa_1
XFILLER_126_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_2_88_2 U$$4306/X U$$4439/X input243/X VGND VGND VPWR VPWR dadda_fa_3_89_1/A
+ dadda_fa_3_88_3/A sky130_fd_sc_hd__fa_1
XFILLER_28_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_956 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdadda_fa_5_65_1 dadda_fa_5_65_1/A dadda_fa_5_65_1/B dadda_fa_5_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_66_0/B dadda_fa_7_65_0/A sky130_fd_sc_hd__fa_1
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_58_0 dadda_fa_5_58_0/A dadda_fa_5_58_0/B dadda_fa_5_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_59_0/A dadda_fa_6_58_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
.ends

