VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Microwatt_FP_DFFRFile
  CLASS BLOCK ;
  FOREIGN Microwatt_FP_DFFRFile ;
  ORIGIN 0.000 0.000 ;
  SIZE 1150.000 BY 1150.000 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 1146.000 21.530 1150.000 ;
    END
  END CLK
  PIN D1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END D1[0]
  PIN D1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END D1[10]
  PIN D1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END D1[11]
  PIN D1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END D1[12]
  PIN D1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END D1[13]
  PIN D1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END D1[14]
  PIN D1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END D1[15]
  PIN D1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END D1[16]
  PIN D1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END D1[17]
  PIN D1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END D1[18]
  PIN D1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END D1[19]
  PIN D1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END D1[1]
  PIN D1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END D1[20]
  PIN D1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END D1[21]
  PIN D1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END D1[22]
  PIN D1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END D1[23]
  PIN D1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END D1[24]
  PIN D1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END D1[25]
  PIN D1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END D1[26]
  PIN D1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END D1[27]
  PIN D1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END D1[28]
  PIN D1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END D1[29]
  PIN D1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END D1[2]
  PIN D1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END D1[30]
  PIN D1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END D1[31]
  PIN D1[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END D1[32]
  PIN D1[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END D1[33]
  PIN D1[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.520 4.000 314.120 ;
    END
  END D1[34]
  PIN D1[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END D1[35]
  PIN D1[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END D1[36]
  PIN D1[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END D1[37]
  PIN D1[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END D1[38]
  PIN D1[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END D1[39]
  PIN D1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END D1[3]
  PIN D1[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END D1[40]
  PIN D1[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END D1[41]
  PIN D1[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END D1[42]
  PIN D1[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END D1[43]
  PIN D1[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END D1[44]
  PIN D1[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END D1[45]
  PIN D1[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 419.600 4.000 420.200 ;
    END
  END D1[46]
  PIN D1[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END D1[47]
  PIN D1[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.280 4.000 437.880 ;
    END
  END D1[48]
  PIN D1[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END D1[49]
  PIN D1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END D1[4]
  PIN D1[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.960 4.000 455.560 ;
    END
  END D1[50]
  PIN D1[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END D1[51]
  PIN D1[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END D1[52]
  PIN D1[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END D1[53]
  PIN D1[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 490.320 4.000 490.920 ;
    END
  END D1[54]
  PIN D1[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END D1[55]
  PIN D1[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.000 4.000 508.600 ;
    END
  END D1[56]
  PIN D1[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END D1[57]
  PIN D1[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.680 4.000 526.280 ;
    END
  END D1[58]
  PIN D1[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END D1[59]
  PIN D1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END D1[5]
  PIN D1[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END D1[60]
  PIN D1[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END D1[61]
  PIN D1[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END D1[62]
  PIN D1[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END D1[63]
  PIN D1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END D1[6]
  PIN D1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END D1[7]
  PIN D1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END D1[8]
  PIN D1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END D1[9]
  PIN D2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END D2[0]
  PIN D2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.120 4.000 667.720 ;
    END
  END D2[10]
  PIN D2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END D2[11]
  PIN D2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.800 4.000 685.400 ;
    END
  END D2[12]
  PIN D2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END D2[13]
  PIN D2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 702.480 4.000 703.080 ;
    END
  END D2[14]
  PIN D2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 711.320 4.000 711.920 ;
    END
  END D2[15]
  PIN D2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.160 4.000 720.760 ;
    END
  END D2[16]
  PIN D2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.000 4.000 729.600 ;
    END
  END D2[17]
  PIN D2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END D2[18]
  PIN D2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END D2[19]
  PIN D2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END D2[1]
  PIN D2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 755.520 4.000 756.120 ;
    END
  END D2[20]
  PIN D2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 764.360 4.000 764.960 ;
    END
  END D2[21]
  PIN D2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.200 4.000 773.800 ;
    END
  END D2[22]
  PIN D2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END D2[23]
  PIN D2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 790.880 4.000 791.480 ;
    END
  END D2[24]
  PIN D2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.720 4.000 800.320 ;
    END
  END D2[25]
  PIN D2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 808.560 4.000 809.160 ;
    END
  END D2[26]
  PIN D2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END D2[27]
  PIN D2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END D2[28]
  PIN D2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.080 4.000 835.680 ;
    END
  END D2[29]
  PIN D2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 596.400 4.000 597.000 ;
    END
  END D2[2]
  PIN D2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.920 4.000 844.520 ;
    END
  END D2[30]
  PIN D2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 852.760 4.000 853.360 ;
    END
  END D2[31]
  PIN D2[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 861.600 4.000 862.200 ;
    END
  END D2[32]
  PIN D2[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END D2[33]
  PIN D2[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 879.280 4.000 879.880 ;
    END
  END D2[34]
  PIN D2[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END D2[35]
  PIN D2[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.960 4.000 897.560 ;
    END
  END D2[36]
  PIN D2[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.800 4.000 906.400 ;
    END
  END D2[37]
  PIN D2[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 914.640 4.000 915.240 ;
    END
  END D2[38]
  PIN D2[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 923.480 4.000 924.080 ;
    END
  END D2[39]
  PIN D2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END D2[3]
  PIN D2[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 932.320 4.000 932.920 ;
    END
  END D2[40]
  PIN D2[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.160 4.000 941.760 ;
    END
  END D2[41]
  PIN D2[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.000 4.000 950.600 ;
    END
  END D2[42]
  PIN D2[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END D2[43]
  PIN D2[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 967.680 4.000 968.280 ;
    END
  END D2[44]
  PIN D2[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 976.520 4.000 977.120 ;
    END
  END D2[45]
  PIN D2[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 985.360 4.000 985.960 ;
    END
  END D2[46]
  PIN D2[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.200 4.000 994.800 ;
    END
  END D2[47]
  PIN D2[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END D2[48]
  PIN D2[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.880 4.000 1012.480 ;
    END
  END D2[49]
  PIN D2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.080 4.000 614.680 ;
    END
  END D2[4]
  PIN D2[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.720 4.000 1021.320 ;
    END
  END D2[50]
  PIN D2[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1029.560 4.000 1030.160 ;
    END
  END D2[51]
  PIN D2[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1038.400 4.000 1039.000 ;
    END
  END D2[52]
  PIN D2[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END D2[53]
  PIN D2[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.080 4.000 1056.680 ;
    END
  END D2[54]
  PIN D2[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.920 4.000 1065.520 ;
    END
  END D2[55]
  PIN D2[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1073.760 4.000 1074.360 ;
    END
  END D2[56]
  PIN D2[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1082.600 4.000 1083.200 ;
    END
  END D2[57]
  PIN D2[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END D2[58]
  PIN D2[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1100.280 4.000 1100.880 ;
    END
  END D2[59]
  PIN D2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END D2[5]
  PIN D2[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1109.120 4.000 1109.720 ;
    END
  END D2[60]
  PIN D2[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1117.960 4.000 1118.560 ;
    END
  END D2[61]
  PIN D2[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1126.800 4.000 1127.400 ;
    END
  END D2[62]
  PIN D2[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1135.640 4.000 1136.240 ;
    END
  END D2[63]
  PIN D2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END D2[6]
  PIN D2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END D2[7]
  PIN D2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END D2[8]
  PIN D2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END D2[9]
  PIN D3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END D3[0]
  PIN D3[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END D3[10]
  PIN D3[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END D3[11]
  PIN D3[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END D3[12]
  PIN D3[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END D3[13]
  PIN D3[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END D3[14]
  PIN D3[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END D3[15]
  PIN D3[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END D3[16]
  PIN D3[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END D3[17]
  PIN D3[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END D3[18]
  PIN D3[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END D3[19]
  PIN D3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END D3[1]
  PIN D3[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END D3[20]
  PIN D3[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END D3[21]
  PIN D3[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END D3[22]
  PIN D3[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END D3[23]
  PIN D3[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END D3[24]
  PIN D3[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END D3[25]
  PIN D3[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END D3[26]
  PIN D3[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END D3[27]
  PIN D3[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END D3[28]
  PIN D3[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END D3[29]
  PIN D3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END D3[2]
  PIN D3[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END D3[30]
  PIN D3[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END D3[31]
  PIN D3[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END D3[32]
  PIN D3[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END D3[33]
  PIN D3[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END D3[34]
  PIN D3[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END D3[35]
  PIN D3[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 0.000 334.790 4.000 ;
    END
  END D3[36]
  PIN D3[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END D3[37]
  PIN D3[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END D3[38]
  PIN D3[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END D3[39]
  PIN D3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END D3[3]
  PIN D3[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END D3[40]
  PIN D3[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END D3[41]
  PIN D3[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END D3[42]
  PIN D3[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END D3[43]
  PIN D3[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END D3[44]
  PIN D3[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END D3[45]
  PIN D3[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END D3[46]
  PIN D3[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END D3[47]
  PIN D3[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END D3[48]
  PIN D3[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 0.000 448.410 4.000 ;
    END
  END D3[49]
  PIN D3[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END D3[4]
  PIN D3[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 0.000 457.150 4.000 ;
    END
  END D3[50]
  PIN D3[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END D3[51]
  PIN D3[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END D3[52]
  PIN D3[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END D3[53]
  PIN D3[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END D3[54]
  PIN D3[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END D3[55]
  PIN D3[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END D3[56]
  PIN D3[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END D3[57]
  PIN D3[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 0.000 527.070 4.000 ;
    END
  END D3[58]
  PIN D3[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 4.000 ;
    END
  END D3[59]
  PIN D3[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END D3[5]
  PIN D3[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END D3[60]
  PIN D3[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END D3[61]
  PIN D3[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END D3[62]
  PIN D3[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END D3[63]
  PIN D3[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END D3[6]
  PIN D3[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END D3[7]
  PIN D3[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END D3[8]
  PIN D3[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END D3[9]
  PIN DW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 4.000 ;
    END
  END DW[0]
  PIN DW[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END DW[10]
  PIN DW[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 0.000 675.650 4.000 ;
    END
  END DW[11]
  PIN DW[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 4.000 ;
    END
  END DW[12]
  PIN DW[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END DW[13]
  PIN DW[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 0.000 701.870 4.000 ;
    END
  END DW[14]
  PIN DW[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 0.000 710.610 4.000 ;
    END
  END DW[15]
  PIN DW[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 0.000 719.350 4.000 ;
    END
  END DW[16]
  PIN DW[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END DW[17]
  PIN DW[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 0.000 736.830 4.000 ;
    END
  END DW[18]
  PIN DW[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 4.000 ;
    END
  END DW[19]
  PIN DW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END DW[1]
  PIN DW[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 0.000 754.310 4.000 ;
    END
  END DW[20]
  PIN DW[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 0.000 763.050 4.000 ;
    END
  END DW[21]
  PIN DW[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 0.000 771.790 4.000 ;
    END
  END DW[22]
  PIN DW[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END DW[23]
  PIN DW[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END DW[24]
  PIN DW[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END DW[25]
  PIN DW[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 0.000 806.750 4.000 ;
    END
  END DW[26]
  PIN DW[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 0.000 815.490 4.000 ;
    END
  END DW[27]
  PIN DW[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 0.000 824.230 4.000 ;
    END
  END DW[28]
  PIN DW[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 0.000 832.970 4.000 ;
    END
  END DW[29]
  PIN DW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 4.000 ;
    END
  END DW[2]
  PIN DW[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.430 0.000 841.710 4.000 ;
    END
  END DW[30]
  PIN DW[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 0.000 850.450 4.000 ;
    END
  END DW[31]
  PIN DW[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.910 0.000 859.190 4.000 ;
    END
  END DW[32]
  PIN DW[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.650 0.000 867.930 4.000 ;
    END
  END DW[33]
  PIN DW[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 0.000 876.670 4.000 ;
    END
  END DW[34]
  PIN DW[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 0.000 885.410 4.000 ;
    END
  END DW[35]
  PIN DW[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 0.000 894.150 4.000 ;
    END
  END DW[36]
  PIN DW[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 0.000 902.890 4.000 ;
    END
  END DW[37]
  PIN DW[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END DW[38]
  PIN DW[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090 0.000 920.370 4.000 ;
    END
  END DW[39]
  PIN DW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END DW[3]
  PIN DW[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.830 0.000 929.110 4.000 ;
    END
  END DW[40]
  PIN DW[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.570 0.000 937.850 4.000 ;
    END
  END DW[41]
  PIN DW[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 0.000 946.590 4.000 ;
    END
  END DW[42]
  PIN DW[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 0.000 955.330 4.000 ;
    END
  END DW[43]
  PIN DW[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.790 0.000 964.070 4.000 ;
    END
  END DW[44]
  PIN DW[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END DW[45]
  PIN DW[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 0.000 981.550 4.000 ;
    END
  END DW[46]
  PIN DW[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 0.000 990.290 4.000 ;
    END
  END DW[47]
  PIN DW[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 0.000 999.030 4.000 ;
    END
  END DW[48]
  PIN DW[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.490 0.000 1007.770 4.000 ;
    END
  END DW[49]
  PIN DW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END DW[4]
  PIN DW[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.230 0.000 1016.510 4.000 ;
    END
  END DW[50]
  PIN DW[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.970 0.000 1025.250 4.000 ;
    END
  END DW[51]
  PIN DW[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END DW[52]
  PIN DW[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.450 0.000 1042.730 4.000 ;
    END
  END DW[53]
  PIN DW[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 0.000 1051.470 4.000 ;
    END
  END DW[54]
  PIN DW[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.930 0.000 1060.210 4.000 ;
    END
  END DW[55]
  PIN DW[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.670 0.000 1068.950 4.000 ;
    END
  END DW[56]
  PIN DW[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.410 0.000 1077.690 4.000 ;
    END
  END DW[57]
  PIN DW[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.150 0.000 1086.430 4.000 ;
    END
  END DW[58]
  PIN DW[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END DW[59]
  PIN DW[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END DW[5]
  PIN DW[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.630 0.000 1103.910 4.000 ;
    END
  END DW[60]
  PIN DW[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.370 0.000 1112.650 4.000 ;
    END
  END DW[61]
  PIN DW[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 0.000 1121.390 4.000 ;
    END
  END DW[62]
  PIN DW[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.850 0.000 1130.130 4.000 ;
    END
  END DW[63]
  PIN DW[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 0.000 631.950 4.000 ;
    END
  END DW[6]
  PIN DW[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END DW[7]
  PIN DW[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 4.000 ;
    END
  END DW[8]
  PIN DW[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END DW[9]
  PIN R1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 1146.000 97.890 1150.000 ;
    END
  END R1[0]
  PIN R1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 1146.000 136.070 1150.000 ;
    END
  END R1[1]
  PIN R1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 1146.000 174.250 1150.000 ;
    END
  END R1[2]
  PIN R1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 1146.000 212.430 1150.000 ;
    END
  END R1[3]
  PIN R1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 1146.000 250.610 1150.000 ;
    END
  END R1[4]
  PIN R1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 1146.000 288.790 1150.000 ;
    END
  END R1[5]
  PIN R1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 1146.000 326.970 1150.000 ;
    END
  END R1[6]
  PIN R2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 1146.000 365.150 1150.000 ;
    END
  END R2[0]
  PIN R2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 1146.000 403.330 1150.000 ;
    END
  END R2[1]
  PIN R2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 1146.000 441.510 1150.000 ;
    END
  END R2[2]
  PIN R2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 1146.000 479.690 1150.000 ;
    END
  END R2[3]
  PIN R2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 1146.000 517.870 1150.000 ;
    END
  END R2[4]
  PIN R2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 1146.000 556.050 1150.000 ;
    END
  END R2[5]
  PIN R2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 1146.000 594.230 1150.000 ;
    END
  END R2[6]
  PIN R3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 1146.000 632.410 1150.000 ;
    END
  END R3[0]
  PIN R3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 1146.000 670.590 1150.000 ;
    END
  END R3[1]
  PIN R3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 1146.000 708.770 1150.000 ;
    END
  END R3[2]
  PIN R3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 1146.000 746.950 1150.000 ;
    END
  END R3[3]
  PIN R3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 1146.000 785.130 1150.000 ;
    END
  END R3[4]
  PIN R3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.030 1146.000 823.310 1150.000 ;
    END
  END R3[5]
  PIN R3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 1146.000 861.490 1150.000 ;
    END
  END R3[6]
  PIN RW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 1146.000 899.670 1150.000 ;
    END
  END RW[0]
  PIN RW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.570 1146.000 937.850 1150.000 ;
    END
  END RW[1]
  PIN RW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 1146.000 976.030 1150.000 ;
    END
  END RW[2]
  PIN RW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.930 1146.000 1014.210 1150.000 ;
    END
  END RW[3]
  PIN RW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.110 1146.000 1052.390 1150.000 ;
    END
  END RW[4]
  PIN RW[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.290 1146.000 1090.570 1150.000 ;
    END
  END RW[5]
  PIN RW[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.470 1146.000 1128.750 1150.000 ;
    END
  END RW[6]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 98.970 10.640 102.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 10.640 282.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 10.640 462.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 10.640 642.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 10.640 822.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 10.640 1002.070 1137.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.970 10.640 12.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 10.640 192.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 10.640 372.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 10.640 552.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 10.640 732.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 10.640 912.070 1137.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 10.640 1092.070 1137.200 ;
    END
  END VPWR
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 1146.000 59.710 1150.000 ;
    END
  END WE
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1144.480 1137.045 ;
      LAYER met1 ;
        RECT 2.830 2.420 1144.480 1137.200 ;
      LAYER met2 ;
        RECT 2.860 1145.720 20.970 1146.000 ;
        RECT 21.810 1145.720 59.150 1146.000 ;
        RECT 59.990 1145.720 97.330 1146.000 ;
        RECT 98.170 1145.720 135.510 1146.000 ;
        RECT 136.350 1145.720 173.690 1146.000 ;
        RECT 174.530 1145.720 211.870 1146.000 ;
        RECT 212.710 1145.720 250.050 1146.000 ;
        RECT 250.890 1145.720 288.230 1146.000 ;
        RECT 289.070 1145.720 326.410 1146.000 ;
        RECT 327.250 1145.720 364.590 1146.000 ;
        RECT 365.430 1145.720 402.770 1146.000 ;
        RECT 403.610 1145.720 440.950 1146.000 ;
        RECT 441.790 1145.720 479.130 1146.000 ;
        RECT 479.970 1145.720 517.310 1146.000 ;
        RECT 518.150 1145.720 555.490 1146.000 ;
        RECT 556.330 1145.720 593.670 1146.000 ;
        RECT 594.510 1145.720 631.850 1146.000 ;
        RECT 632.690 1145.720 670.030 1146.000 ;
        RECT 670.870 1145.720 708.210 1146.000 ;
        RECT 709.050 1145.720 746.390 1146.000 ;
        RECT 747.230 1145.720 784.570 1146.000 ;
        RECT 785.410 1145.720 822.750 1146.000 ;
        RECT 823.590 1145.720 860.930 1146.000 ;
        RECT 861.770 1145.720 899.110 1146.000 ;
        RECT 899.950 1145.720 937.290 1146.000 ;
        RECT 938.130 1145.720 975.470 1146.000 ;
        RECT 976.310 1145.720 1013.650 1146.000 ;
        RECT 1014.490 1145.720 1051.830 1146.000 ;
        RECT 1052.670 1145.720 1090.010 1146.000 ;
        RECT 1090.850 1145.720 1128.190 1146.000 ;
        RECT 1129.030 1145.720 1141.160 1146.000 ;
        RECT 2.860 4.280 1141.160 1145.720 ;
        RECT 2.860 2.390 19.590 4.280 ;
        RECT 20.430 2.390 28.330 4.280 ;
        RECT 29.170 2.390 37.070 4.280 ;
        RECT 37.910 2.390 45.810 4.280 ;
        RECT 46.650 2.390 54.550 4.280 ;
        RECT 55.390 2.390 63.290 4.280 ;
        RECT 64.130 2.390 72.030 4.280 ;
        RECT 72.870 2.390 80.770 4.280 ;
        RECT 81.610 2.390 89.510 4.280 ;
        RECT 90.350 2.390 98.250 4.280 ;
        RECT 99.090 2.390 106.990 4.280 ;
        RECT 107.830 2.390 115.730 4.280 ;
        RECT 116.570 2.390 124.470 4.280 ;
        RECT 125.310 2.390 133.210 4.280 ;
        RECT 134.050 2.390 141.950 4.280 ;
        RECT 142.790 2.390 150.690 4.280 ;
        RECT 151.530 2.390 159.430 4.280 ;
        RECT 160.270 2.390 168.170 4.280 ;
        RECT 169.010 2.390 176.910 4.280 ;
        RECT 177.750 2.390 185.650 4.280 ;
        RECT 186.490 2.390 194.390 4.280 ;
        RECT 195.230 2.390 203.130 4.280 ;
        RECT 203.970 2.390 211.870 4.280 ;
        RECT 212.710 2.390 220.610 4.280 ;
        RECT 221.450 2.390 229.350 4.280 ;
        RECT 230.190 2.390 238.090 4.280 ;
        RECT 238.930 2.390 246.830 4.280 ;
        RECT 247.670 2.390 255.570 4.280 ;
        RECT 256.410 2.390 264.310 4.280 ;
        RECT 265.150 2.390 273.050 4.280 ;
        RECT 273.890 2.390 281.790 4.280 ;
        RECT 282.630 2.390 290.530 4.280 ;
        RECT 291.370 2.390 299.270 4.280 ;
        RECT 300.110 2.390 308.010 4.280 ;
        RECT 308.850 2.390 316.750 4.280 ;
        RECT 317.590 2.390 325.490 4.280 ;
        RECT 326.330 2.390 334.230 4.280 ;
        RECT 335.070 2.390 342.970 4.280 ;
        RECT 343.810 2.390 351.710 4.280 ;
        RECT 352.550 2.390 360.450 4.280 ;
        RECT 361.290 2.390 369.190 4.280 ;
        RECT 370.030 2.390 377.930 4.280 ;
        RECT 378.770 2.390 386.670 4.280 ;
        RECT 387.510 2.390 395.410 4.280 ;
        RECT 396.250 2.390 404.150 4.280 ;
        RECT 404.990 2.390 412.890 4.280 ;
        RECT 413.730 2.390 421.630 4.280 ;
        RECT 422.470 2.390 430.370 4.280 ;
        RECT 431.210 2.390 439.110 4.280 ;
        RECT 439.950 2.390 447.850 4.280 ;
        RECT 448.690 2.390 456.590 4.280 ;
        RECT 457.430 2.390 465.330 4.280 ;
        RECT 466.170 2.390 474.070 4.280 ;
        RECT 474.910 2.390 482.810 4.280 ;
        RECT 483.650 2.390 491.550 4.280 ;
        RECT 492.390 2.390 500.290 4.280 ;
        RECT 501.130 2.390 509.030 4.280 ;
        RECT 509.870 2.390 517.770 4.280 ;
        RECT 518.610 2.390 526.510 4.280 ;
        RECT 527.350 2.390 535.250 4.280 ;
        RECT 536.090 2.390 543.990 4.280 ;
        RECT 544.830 2.390 552.730 4.280 ;
        RECT 553.570 2.390 561.470 4.280 ;
        RECT 562.310 2.390 570.210 4.280 ;
        RECT 571.050 2.390 578.950 4.280 ;
        RECT 579.790 2.390 587.690 4.280 ;
        RECT 588.530 2.390 596.430 4.280 ;
        RECT 597.270 2.390 605.170 4.280 ;
        RECT 606.010 2.390 613.910 4.280 ;
        RECT 614.750 2.390 622.650 4.280 ;
        RECT 623.490 2.390 631.390 4.280 ;
        RECT 632.230 2.390 640.130 4.280 ;
        RECT 640.970 2.390 648.870 4.280 ;
        RECT 649.710 2.390 657.610 4.280 ;
        RECT 658.450 2.390 666.350 4.280 ;
        RECT 667.190 2.390 675.090 4.280 ;
        RECT 675.930 2.390 683.830 4.280 ;
        RECT 684.670 2.390 692.570 4.280 ;
        RECT 693.410 2.390 701.310 4.280 ;
        RECT 702.150 2.390 710.050 4.280 ;
        RECT 710.890 2.390 718.790 4.280 ;
        RECT 719.630 2.390 727.530 4.280 ;
        RECT 728.370 2.390 736.270 4.280 ;
        RECT 737.110 2.390 745.010 4.280 ;
        RECT 745.850 2.390 753.750 4.280 ;
        RECT 754.590 2.390 762.490 4.280 ;
        RECT 763.330 2.390 771.230 4.280 ;
        RECT 772.070 2.390 779.970 4.280 ;
        RECT 780.810 2.390 788.710 4.280 ;
        RECT 789.550 2.390 797.450 4.280 ;
        RECT 798.290 2.390 806.190 4.280 ;
        RECT 807.030 2.390 814.930 4.280 ;
        RECT 815.770 2.390 823.670 4.280 ;
        RECT 824.510 2.390 832.410 4.280 ;
        RECT 833.250 2.390 841.150 4.280 ;
        RECT 841.990 2.390 849.890 4.280 ;
        RECT 850.730 2.390 858.630 4.280 ;
        RECT 859.470 2.390 867.370 4.280 ;
        RECT 868.210 2.390 876.110 4.280 ;
        RECT 876.950 2.390 884.850 4.280 ;
        RECT 885.690 2.390 893.590 4.280 ;
        RECT 894.430 2.390 902.330 4.280 ;
        RECT 903.170 2.390 911.070 4.280 ;
        RECT 911.910 2.390 919.810 4.280 ;
        RECT 920.650 2.390 928.550 4.280 ;
        RECT 929.390 2.390 937.290 4.280 ;
        RECT 938.130 2.390 946.030 4.280 ;
        RECT 946.870 2.390 954.770 4.280 ;
        RECT 955.610 2.390 963.510 4.280 ;
        RECT 964.350 2.390 972.250 4.280 ;
        RECT 973.090 2.390 980.990 4.280 ;
        RECT 981.830 2.390 989.730 4.280 ;
        RECT 990.570 2.390 998.470 4.280 ;
        RECT 999.310 2.390 1007.210 4.280 ;
        RECT 1008.050 2.390 1015.950 4.280 ;
        RECT 1016.790 2.390 1024.690 4.280 ;
        RECT 1025.530 2.390 1033.430 4.280 ;
        RECT 1034.270 2.390 1042.170 4.280 ;
        RECT 1043.010 2.390 1050.910 4.280 ;
        RECT 1051.750 2.390 1059.650 4.280 ;
        RECT 1060.490 2.390 1068.390 4.280 ;
        RECT 1069.230 2.390 1077.130 4.280 ;
        RECT 1077.970 2.390 1085.870 4.280 ;
        RECT 1086.710 2.390 1094.610 4.280 ;
        RECT 1095.450 2.390 1103.350 4.280 ;
        RECT 1104.190 2.390 1112.090 4.280 ;
        RECT 1112.930 2.390 1120.830 4.280 ;
        RECT 1121.670 2.390 1129.570 4.280 ;
        RECT 1130.410 2.390 1141.160 4.280 ;
      LAYER met3 ;
        RECT 3.745 1136.640 1136.595 1137.125 ;
        RECT 4.400 1135.240 1136.595 1136.640 ;
        RECT 3.745 1127.800 1136.595 1135.240 ;
        RECT 4.400 1126.400 1136.595 1127.800 ;
        RECT 3.745 1118.960 1136.595 1126.400 ;
        RECT 4.400 1117.560 1136.595 1118.960 ;
        RECT 3.745 1110.120 1136.595 1117.560 ;
        RECT 4.400 1108.720 1136.595 1110.120 ;
        RECT 3.745 1101.280 1136.595 1108.720 ;
        RECT 4.400 1099.880 1136.595 1101.280 ;
        RECT 3.745 1092.440 1136.595 1099.880 ;
        RECT 4.400 1091.040 1136.595 1092.440 ;
        RECT 3.745 1083.600 1136.595 1091.040 ;
        RECT 4.400 1082.200 1136.595 1083.600 ;
        RECT 3.745 1074.760 1136.595 1082.200 ;
        RECT 4.400 1073.360 1136.595 1074.760 ;
        RECT 3.745 1065.920 1136.595 1073.360 ;
        RECT 4.400 1064.520 1136.595 1065.920 ;
        RECT 3.745 1057.080 1136.595 1064.520 ;
        RECT 4.400 1055.680 1136.595 1057.080 ;
        RECT 3.745 1048.240 1136.595 1055.680 ;
        RECT 4.400 1046.840 1136.595 1048.240 ;
        RECT 3.745 1039.400 1136.595 1046.840 ;
        RECT 4.400 1038.000 1136.595 1039.400 ;
        RECT 3.745 1030.560 1136.595 1038.000 ;
        RECT 4.400 1029.160 1136.595 1030.560 ;
        RECT 3.745 1021.720 1136.595 1029.160 ;
        RECT 4.400 1020.320 1136.595 1021.720 ;
        RECT 3.745 1012.880 1136.595 1020.320 ;
        RECT 4.400 1011.480 1136.595 1012.880 ;
        RECT 3.745 1004.040 1136.595 1011.480 ;
        RECT 4.400 1002.640 1136.595 1004.040 ;
        RECT 3.745 995.200 1136.595 1002.640 ;
        RECT 4.400 993.800 1136.595 995.200 ;
        RECT 3.745 986.360 1136.595 993.800 ;
        RECT 4.400 984.960 1136.595 986.360 ;
        RECT 3.745 977.520 1136.595 984.960 ;
        RECT 4.400 976.120 1136.595 977.520 ;
        RECT 3.745 968.680 1136.595 976.120 ;
        RECT 4.400 967.280 1136.595 968.680 ;
        RECT 3.745 959.840 1136.595 967.280 ;
        RECT 4.400 958.440 1136.595 959.840 ;
        RECT 3.745 951.000 1136.595 958.440 ;
        RECT 4.400 949.600 1136.595 951.000 ;
        RECT 3.745 942.160 1136.595 949.600 ;
        RECT 4.400 940.760 1136.595 942.160 ;
        RECT 3.745 933.320 1136.595 940.760 ;
        RECT 4.400 931.920 1136.595 933.320 ;
        RECT 3.745 924.480 1136.595 931.920 ;
        RECT 4.400 923.080 1136.595 924.480 ;
        RECT 3.745 915.640 1136.595 923.080 ;
        RECT 4.400 914.240 1136.595 915.640 ;
        RECT 3.745 906.800 1136.595 914.240 ;
        RECT 4.400 905.400 1136.595 906.800 ;
        RECT 3.745 897.960 1136.595 905.400 ;
        RECT 4.400 896.560 1136.595 897.960 ;
        RECT 3.745 889.120 1136.595 896.560 ;
        RECT 4.400 887.720 1136.595 889.120 ;
        RECT 3.745 880.280 1136.595 887.720 ;
        RECT 4.400 878.880 1136.595 880.280 ;
        RECT 3.745 871.440 1136.595 878.880 ;
        RECT 4.400 870.040 1136.595 871.440 ;
        RECT 3.745 862.600 1136.595 870.040 ;
        RECT 4.400 861.200 1136.595 862.600 ;
        RECT 3.745 853.760 1136.595 861.200 ;
        RECT 4.400 852.360 1136.595 853.760 ;
        RECT 3.745 844.920 1136.595 852.360 ;
        RECT 4.400 843.520 1136.595 844.920 ;
        RECT 3.745 836.080 1136.595 843.520 ;
        RECT 4.400 834.680 1136.595 836.080 ;
        RECT 3.745 827.240 1136.595 834.680 ;
        RECT 4.400 825.840 1136.595 827.240 ;
        RECT 3.745 818.400 1136.595 825.840 ;
        RECT 4.400 817.000 1136.595 818.400 ;
        RECT 3.745 809.560 1136.595 817.000 ;
        RECT 4.400 808.160 1136.595 809.560 ;
        RECT 3.745 800.720 1136.595 808.160 ;
        RECT 4.400 799.320 1136.595 800.720 ;
        RECT 3.745 791.880 1136.595 799.320 ;
        RECT 4.400 790.480 1136.595 791.880 ;
        RECT 3.745 783.040 1136.595 790.480 ;
        RECT 4.400 781.640 1136.595 783.040 ;
        RECT 3.745 774.200 1136.595 781.640 ;
        RECT 4.400 772.800 1136.595 774.200 ;
        RECT 3.745 765.360 1136.595 772.800 ;
        RECT 4.400 763.960 1136.595 765.360 ;
        RECT 3.745 756.520 1136.595 763.960 ;
        RECT 4.400 755.120 1136.595 756.520 ;
        RECT 3.745 747.680 1136.595 755.120 ;
        RECT 4.400 746.280 1136.595 747.680 ;
        RECT 3.745 738.840 1136.595 746.280 ;
        RECT 4.400 737.440 1136.595 738.840 ;
        RECT 3.745 730.000 1136.595 737.440 ;
        RECT 4.400 728.600 1136.595 730.000 ;
        RECT 3.745 721.160 1136.595 728.600 ;
        RECT 4.400 719.760 1136.595 721.160 ;
        RECT 3.745 712.320 1136.595 719.760 ;
        RECT 4.400 710.920 1136.595 712.320 ;
        RECT 3.745 703.480 1136.595 710.920 ;
        RECT 4.400 702.080 1136.595 703.480 ;
        RECT 3.745 694.640 1136.595 702.080 ;
        RECT 4.400 693.240 1136.595 694.640 ;
        RECT 3.745 685.800 1136.595 693.240 ;
        RECT 4.400 684.400 1136.595 685.800 ;
        RECT 3.745 676.960 1136.595 684.400 ;
        RECT 4.400 675.560 1136.595 676.960 ;
        RECT 3.745 668.120 1136.595 675.560 ;
        RECT 4.400 666.720 1136.595 668.120 ;
        RECT 3.745 659.280 1136.595 666.720 ;
        RECT 4.400 657.880 1136.595 659.280 ;
        RECT 3.745 650.440 1136.595 657.880 ;
        RECT 4.400 649.040 1136.595 650.440 ;
        RECT 3.745 641.600 1136.595 649.040 ;
        RECT 4.400 640.200 1136.595 641.600 ;
        RECT 3.745 632.760 1136.595 640.200 ;
        RECT 4.400 631.360 1136.595 632.760 ;
        RECT 3.745 623.920 1136.595 631.360 ;
        RECT 4.400 622.520 1136.595 623.920 ;
        RECT 3.745 615.080 1136.595 622.520 ;
        RECT 4.400 613.680 1136.595 615.080 ;
        RECT 3.745 606.240 1136.595 613.680 ;
        RECT 4.400 604.840 1136.595 606.240 ;
        RECT 3.745 597.400 1136.595 604.840 ;
        RECT 4.400 596.000 1136.595 597.400 ;
        RECT 3.745 588.560 1136.595 596.000 ;
        RECT 4.400 587.160 1136.595 588.560 ;
        RECT 3.745 579.720 1136.595 587.160 ;
        RECT 4.400 578.320 1136.595 579.720 ;
        RECT 3.745 570.880 1136.595 578.320 ;
        RECT 4.400 569.480 1136.595 570.880 ;
        RECT 3.745 562.040 1136.595 569.480 ;
        RECT 4.400 560.640 1136.595 562.040 ;
        RECT 3.745 553.200 1136.595 560.640 ;
        RECT 4.400 551.800 1136.595 553.200 ;
        RECT 3.745 544.360 1136.595 551.800 ;
        RECT 4.400 542.960 1136.595 544.360 ;
        RECT 3.745 535.520 1136.595 542.960 ;
        RECT 4.400 534.120 1136.595 535.520 ;
        RECT 3.745 526.680 1136.595 534.120 ;
        RECT 4.400 525.280 1136.595 526.680 ;
        RECT 3.745 517.840 1136.595 525.280 ;
        RECT 4.400 516.440 1136.595 517.840 ;
        RECT 3.745 509.000 1136.595 516.440 ;
        RECT 4.400 507.600 1136.595 509.000 ;
        RECT 3.745 500.160 1136.595 507.600 ;
        RECT 4.400 498.760 1136.595 500.160 ;
        RECT 3.745 491.320 1136.595 498.760 ;
        RECT 4.400 489.920 1136.595 491.320 ;
        RECT 3.745 482.480 1136.595 489.920 ;
        RECT 4.400 481.080 1136.595 482.480 ;
        RECT 3.745 473.640 1136.595 481.080 ;
        RECT 4.400 472.240 1136.595 473.640 ;
        RECT 3.745 464.800 1136.595 472.240 ;
        RECT 4.400 463.400 1136.595 464.800 ;
        RECT 3.745 455.960 1136.595 463.400 ;
        RECT 4.400 454.560 1136.595 455.960 ;
        RECT 3.745 447.120 1136.595 454.560 ;
        RECT 4.400 445.720 1136.595 447.120 ;
        RECT 3.745 438.280 1136.595 445.720 ;
        RECT 4.400 436.880 1136.595 438.280 ;
        RECT 3.745 429.440 1136.595 436.880 ;
        RECT 4.400 428.040 1136.595 429.440 ;
        RECT 3.745 420.600 1136.595 428.040 ;
        RECT 4.400 419.200 1136.595 420.600 ;
        RECT 3.745 411.760 1136.595 419.200 ;
        RECT 4.400 410.360 1136.595 411.760 ;
        RECT 3.745 402.920 1136.595 410.360 ;
        RECT 4.400 401.520 1136.595 402.920 ;
        RECT 3.745 394.080 1136.595 401.520 ;
        RECT 4.400 392.680 1136.595 394.080 ;
        RECT 3.745 385.240 1136.595 392.680 ;
        RECT 4.400 383.840 1136.595 385.240 ;
        RECT 3.745 376.400 1136.595 383.840 ;
        RECT 4.400 375.000 1136.595 376.400 ;
        RECT 3.745 367.560 1136.595 375.000 ;
        RECT 4.400 366.160 1136.595 367.560 ;
        RECT 3.745 358.720 1136.595 366.160 ;
        RECT 4.400 357.320 1136.595 358.720 ;
        RECT 3.745 349.880 1136.595 357.320 ;
        RECT 4.400 348.480 1136.595 349.880 ;
        RECT 3.745 341.040 1136.595 348.480 ;
        RECT 4.400 339.640 1136.595 341.040 ;
        RECT 3.745 332.200 1136.595 339.640 ;
        RECT 4.400 330.800 1136.595 332.200 ;
        RECT 3.745 323.360 1136.595 330.800 ;
        RECT 4.400 321.960 1136.595 323.360 ;
        RECT 3.745 314.520 1136.595 321.960 ;
        RECT 4.400 313.120 1136.595 314.520 ;
        RECT 3.745 305.680 1136.595 313.120 ;
        RECT 4.400 304.280 1136.595 305.680 ;
        RECT 3.745 296.840 1136.595 304.280 ;
        RECT 4.400 295.440 1136.595 296.840 ;
        RECT 3.745 288.000 1136.595 295.440 ;
        RECT 4.400 286.600 1136.595 288.000 ;
        RECT 3.745 279.160 1136.595 286.600 ;
        RECT 4.400 277.760 1136.595 279.160 ;
        RECT 3.745 270.320 1136.595 277.760 ;
        RECT 4.400 268.920 1136.595 270.320 ;
        RECT 3.745 261.480 1136.595 268.920 ;
        RECT 4.400 260.080 1136.595 261.480 ;
        RECT 3.745 252.640 1136.595 260.080 ;
        RECT 4.400 251.240 1136.595 252.640 ;
        RECT 3.745 243.800 1136.595 251.240 ;
        RECT 4.400 242.400 1136.595 243.800 ;
        RECT 3.745 234.960 1136.595 242.400 ;
        RECT 4.400 233.560 1136.595 234.960 ;
        RECT 3.745 226.120 1136.595 233.560 ;
        RECT 4.400 224.720 1136.595 226.120 ;
        RECT 3.745 217.280 1136.595 224.720 ;
        RECT 4.400 215.880 1136.595 217.280 ;
        RECT 3.745 208.440 1136.595 215.880 ;
        RECT 4.400 207.040 1136.595 208.440 ;
        RECT 3.745 199.600 1136.595 207.040 ;
        RECT 4.400 198.200 1136.595 199.600 ;
        RECT 3.745 190.760 1136.595 198.200 ;
        RECT 4.400 189.360 1136.595 190.760 ;
        RECT 3.745 181.920 1136.595 189.360 ;
        RECT 4.400 180.520 1136.595 181.920 ;
        RECT 3.745 173.080 1136.595 180.520 ;
        RECT 4.400 171.680 1136.595 173.080 ;
        RECT 3.745 164.240 1136.595 171.680 ;
        RECT 4.400 162.840 1136.595 164.240 ;
        RECT 3.745 155.400 1136.595 162.840 ;
        RECT 4.400 154.000 1136.595 155.400 ;
        RECT 3.745 146.560 1136.595 154.000 ;
        RECT 4.400 145.160 1136.595 146.560 ;
        RECT 3.745 137.720 1136.595 145.160 ;
        RECT 4.400 136.320 1136.595 137.720 ;
        RECT 3.745 128.880 1136.595 136.320 ;
        RECT 4.400 127.480 1136.595 128.880 ;
        RECT 3.745 120.040 1136.595 127.480 ;
        RECT 4.400 118.640 1136.595 120.040 ;
        RECT 3.745 111.200 1136.595 118.640 ;
        RECT 4.400 109.800 1136.595 111.200 ;
        RECT 3.745 102.360 1136.595 109.800 ;
        RECT 4.400 100.960 1136.595 102.360 ;
        RECT 3.745 93.520 1136.595 100.960 ;
        RECT 4.400 92.120 1136.595 93.520 ;
        RECT 3.745 84.680 1136.595 92.120 ;
        RECT 4.400 83.280 1136.595 84.680 ;
        RECT 3.745 75.840 1136.595 83.280 ;
        RECT 4.400 74.440 1136.595 75.840 ;
        RECT 3.745 67.000 1136.595 74.440 ;
        RECT 4.400 65.600 1136.595 67.000 ;
        RECT 3.745 58.160 1136.595 65.600 ;
        RECT 4.400 56.760 1136.595 58.160 ;
        RECT 3.745 49.320 1136.595 56.760 ;
        RECT 4.400 47.920 1136.595 49.320 ;
        RECT 3.745 40.480 1136.595 47.920 ;
        RECT 4.400 39.080 1136.595 40.480 ;
        RECT 3.745 31.640 1136.595 39.080 ;
        RECT 4.400 30.240 1136.595 31.640 ;
        RECT 3.745 22.800 1136.595 30.240 ;
        RECT 4.400 21.400 1136.595 22.800 ;
        RECT 3.745 13.960 1136.595 21.400 ;
        RECT 4.400 12.560 1136.595 13.960 ;
        RECT 3.745 6.975 1136.595 12.560 ;
      LAYER met4 ;
        RECT 4.895 19.895 8.570 1136.105 ;
        RECT 12.470 19.895 98.570 1136.105 ;
        RECT 102.470 19.895 188.570 1136.105 ;
        RECT 192.470 19.895 278.570 1136.105 ;
        RECT 282.470 19.895 368.570 1136.105 ;
        RECT 372.470 19.895 458.570 1136.105 ;
        RECT 462.470 19.895 548.570 1136.105 ;
        RECT 552.470 19.895 638.570 1136.105 ;
        RECT 642.470 19.895 728.570 1136.105 ;
        RECT 732.470 19.895 818.570 1136.105 ;
        RECT 822.470 19.895 908.570 1136.105 ;
        RECT 912.470 19.895 998.570 1136.105 ;
        RECT 1002.470 19.895 1088.570 1136.105 ;
        RECT 1092.470 19.895 1121.185 1136.105 ;
  END
END Microwatt_FP_DFFRFile
END LIBRARY

