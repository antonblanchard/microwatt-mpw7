magic
tech sky130A
magscale 1 2
timestamp 1657539830
<< obsli1 >>
rect 1104 2159 118864 117521
<< obsm1 >>
rect 474 1300 119770 117552
<< metal2 >>
rect 570 119200 626 120000
rect 1490 119200 1546 120000
rect 2410 119200 2466 120000
rect 3330 119200 3386 120000
rect 4250 119200 4306 120000
rect 5170 119200 5226 120000
rect 6090 119200 6146 120000
rect 7010 119200 7066 120000
rect 7930 119200 7986 120000
rect 8850 119200 8906 120000
rect 9770 119200 9826 120000
rect 10690 119200 10746 120000
rect 11610 119200 11666 120000
rect 12530 119200 12586 120000
rect 13450 119200 13506 120000
rect 14370 119200 14426 120000
rect 15290 119200 15346 120000
rect 16210 119200 16266 120000
rect 17130 119200 17186 120000
rect 18050 119200 18106 120000
rect 18970 119200 19026 120000
rect 19890 119200 19946 120000
rect 20810 119200 20866 120000
rect 21730 119200 21786 120000
rect 22650 119200 22706 120000
rect 23570 119200 23626 120000
rect 24490 119200 24546 120000
rect 25410 119200 25466 120000
rect 26330 119200 26386 120000
rect 27250 119200 27306 120000
rect 28170 119200 28226 120000
rect 29090 119200 29146 120000
rect 30010 119200 30066 120000
rect 30930 119200 30986 120000
rect 31850 119200 31906 120000
rect 32770 119200 32826 120000
rect 33690 119200 33746 120000
rect 34610 119200 34666 120000
rect 35530 119200 35586 120000
rect 36450 119200 36506 120000
rect 37370 119200 37426 120000
rect 38290 119200 38346 120000
rect 39210 119200 39266 120000
rect 40130 119200 40186 120000
rect 41050 119200 41106 120000
rect 41970 119200 42026 120000
rect 42890 119200 42946 120000
rect 43810 119200 43866 120000
rect 44730 119200 44786 120000
rect 45650 119200 45706 120000
rect 46570 119200 46626 120000
rect 47490 119200 47546 120000
rect 48410 119200 48466 120000
rect 49330 119200 49386 120000
rect 50250 119200 50306 120000
rect 51170 119200 51226 120000
rect 52090 119200 52146 120000
rect 53010 119200 53066 120000
rect 53930 119200 53986 120000
rect 54850 119200 54906 120000
rect 55770 119200 55826 120000
rect 56690 119200 56746 120000
rect 57610 119200 57666 120000
rect 58530 119200 58586 120000
rect 59450 119200 59506 120000
rect 60370 119200 60426 120000
rect 61290 119200 61346 120000
rect 62210 119200 62266 120000
rect 63130 119200 63186 120000
rect 64050 119200 64106 120000
rect 64970 119200 65026 120000
rect 65890 119200 65946 120000
rect 66810 119200 66866 120000
rect 67730 119200 67786 120000
rect 68650 119200 68706 120000
rect 69570 119200 69626 120000
rect 70490 119200 70546 120000
rect 71410 119200 71466 120000
rect 72330 119200 72386 120000
rect 73250 119200 73306 120000
rect 74170 119200 74226 120000
rect 75090 119200 75146 120000
rect 76010 119200 76066 120000
rect 76930 119200 76986 120000
rect 77850 119200 77906 120000
rect 78770 119200 78826 120000
rect 79690 119200 79746 120000
rect 80610 119200 80666 120000
rect 81530 119200 81586 120000
rect 82450 119200 82506 120000
rect 83370 119200 83426 120000
rect 84290 119200 84346 120000
rect 85210 119200 85266 120000
rect 86130 119200 86186 120000
rect 87050 119200 87106 120000
rect 87970 119200 88026 120000
rect 88890 119200 88946 120000
rect 89810 119200 89866 120000
rect 90730 119200 90786 120000
rect 91650 119200 91706 120000
rect 92570 119200 92626 120000
rect 93490 119200 93546 120000
rect 94410 119200 94466 120000
rect 95330 119200 95386 120000
rect 96250 119200 96306 120000
rect 97170 119200 97226 120000
rect 98090 119200 98146 120000
rect 99010 119200 99066 120000
rect 99930 119200 99986 120000
rect 100850 119200 100906 120000
rect 101770 119200 101826 120000
rect 102690 119200 102746 120000
rect 103610 119200 103666 120000
rect 104530 119200 104586 120000
rect 105450 119200 105506 120000
rect 106370 119200 106426 120000
rect 107290 119200 107346 120000
rect 108210 119200 108266 120000
rect 109130 119200 109186 120000
rect 110050 119200 110106 120000
rect 110970 119200 111026 120000
rect 111890 119200 111946 120000
rect 112810 119200 112866 120000
rect 113730 119200 113786 120000
rect 114650 119200 114706 120000
rect 115570 119200 115626 120000
rect 116490 119200 116546 120000
rect 117410 119200 117466 120000
rect 118330 119200 118386 120000
rect 119250 119200 119306 120000
rect 1490 0 1546 800
rect 2410 0 2466 800
rect 3330 0 3386 800
rect 4250 0 4306 800
rect 5170 0 5226 800
rect 6090 0 6146 800
rect 7010 0 7066 800
rect 7930 0 7986 800
rect 8850 0 8906 800
rect 9770 0 9826 800
rect 10690 0 10746 800
rect 11610 0 11666 800
rect 12530 0 12586 800
rect 13450 0 13506 800
rect 14370 0 14426 800
rect 15290 0 15346 800
rect 16210 0 16266 800
rect 17130 0 17186 800
rect 18050 0 18106 800
rect 18970 0 19026 800
rect 19890 0 19946 800
rect 20810 0 20866 800
rect 21730 0 21786 800
rect 22650 0 22706 800
rect 23570 0 23626 800
rect 24490 0 24546 800
rect 25410 0 25466 800
rect 26330 0 26386 800
rect 27250 0 27306 800
rect 28170 0 28226 800
rect 29090 0 29146 800
rect 30010 0 30066 800
rect 30930 0 30986 800
rect 31850 0 31906 800
rect 32770 0 32826 800
rect 33690 0 33746 800
rect 34610 0 34666 800
rect 35530 0 35586 800
rect 36450 0 36506 800
rect 37370 0 37426 800
rect 38290 0 38346 800
rect 39210 0 39266 800
rect 40130 0 40186 800
rect 41050 0 41106 800
rect 41970 0 42026 800
rect 42890 0 42946 800
rect 43810 0 43866 800
rect 44730 0 44786 800
rect 45650 0 45706 800
rect 46570 0 46626 800
rect 47490 0 47546 800
rect 48410 0 48466 800
rect 49330 0 49386 800
rect 50250 0 50306 800
rect 51170 0 51226 800
rect 52090 0 52146 800
rect 53010 0 53066 800
rect 53930 0 53986 800
rect 54850 0 54906 800
rect 55770 0 55826 800
rect 56690 0 56746 800
rect 57610 0 57666 800
rect 58530 0 58586 800
rect 59450 0 59506 800
rect 60370 0 60426 800
rect 61290 0 61346 800
rect 62210 0 62266 800
rect 63130 0 63186 800
rect 64050 0 64106 800
rect 64970 0 65026 800
rect 65890 0 65946 800
rect 66810 0 66866 800
rect 67730 0 67786 800
rect 68650 0 68706 800
rect 69570 0 69626 800
rect 70490 0 70546 800
rect 71410 0 71466 800
rect 72330 0 72386 800
rect 73250 0 73306 800
rect 74170 0 74226 800
rect 75090 0 75146 800
rect 76010 0 76066 800
rect 76930 0 76986 800
rect 77850 0 77906 800
rect 78770 0 78826 800
rect 79690 0 79746 800
rect 80610 0 80666 800
rect 81530 0 81586 800
rect 82450 0 82506 800
rect 83370 0 83426 800
rect 84290 0 84346 800
rect 85210 0 85266 800
rect 86130 0 86186 800
rect 87050 0 87106 800
rect 87970 0 88026 800
rect 88890 0 88946 800
rect 89810 0 89866 800
rect 90730 0 90786 800
rect 91650 0 91706 800
rect 92570 0 92626 800
rect 93490 0 93546 800
rect 94410 0 94466 800
rect 95330 0 95386 800
rect 96250 0 96306 800
rect 97170 0 97226 800
rect 98090 0 98146 800
rect 99010 0 99066 800
rect 99930 0 99986 800
rect 100850 0 100906 800
rect 101770 0 101826 800
rect 102690 0 102746 800
rect 103610 0 103666 800
rect 104530 0 104586 800
rect 105450 0 105506 800
rect 106370 0 106426 800
rect 107290 0 107346 800
rect 108210 0 108266 800
rect 109130 0 109186 800
rect 110050 0 110106 800
rect 110970 0 111026 800
rect 111890 0 111946 800
rect 112810 0 112866 800
rect 113730 0 113786 800
rect 114650 0 114706 800
rect 115570 0 115626 800
rect 116490 0 116546 800
rect 117410 0 117466 800
rect 118330 0 118386 800
<< obsm2 >>
rect 480 119144 514 119354
rect 682 119144 1434 119354
rect 1602 119144 2354 119354
rect 2522 119144 3274 119354
rect 3442 119144 4194 119354
rect 4362 119144 5114 119354
rect 5282 119144 6034 119354
rect 6202 119144 6954 119354
rect 7122 119144 7874 119354
rect 8042 119144 8794 119354
rect 8962 119144 9714 119354
rect 9882 119144 10634 119354
rect 10802 119144 11554 119354
rect 11722 119144 12474 119354
rect 12642 119144 13394 119354
rect 13562 119144 14314 119354
rect 14482 119144 15234 119354
rect 15402 119144 16154 119354
rect 16322 119144 17074 119354
rect 17242 119144 17994 119354
rect 18162 119144 18914 119354
rect 19082 119144 19834 119354
rect 20002 119144 20754 119354
rect 20922 119144 21674 119354
rect 21842 119144 22594 119354
rect 22762 119144 23514 119354
rect 23682 119144 24434 119354
rect 24602 119144 25354 119354
rect 25522 119144 26274 119354
rect 26442 119144 27194 119354
rect 27362 119144 28114 119354
rect 28282 119144 29034 119354
rect 29202 119144 29954 119354
rect 30122 119144 30874 119354
rect 31042 119144 31794 119354
rect 31962 119144 32714 119354
rect 32882 119144 33634 119354
rect 33802 119144 34554 119354
rect 34722 119144 35474 119354
rect 35642 119144 36394 119354
rect 36562 119144 37314 119354
rect 37482 119144 38234 119354
rect 38402 119144 39154 119354
rect 39322 119144 40074 119354
rect 40242 119144 40994 119354
rect 41162 119144 41914 119354
rect 42082 119144 42834 119354
rect 43002 119144 43754 119354
rect 43922 119144 44674 119354
rect 44842 119144 45594 119354
rect 45762 119144 46514 119354
rect 46682 119144 47434 119354
rect 47602 119144 48354 119354
rect 48522 119144 49274 119354
rect 49442 119144 50194 119354
rect 50362 119144 51114 119354
rect 51282 119144 52034 119354
rect 52202 119144 52954 119354
rect 53122 119144 53874 119354
rect 54042 119144 54794 119354
rect 54962 119144 55714 119354
rect 55882 119144 56634 119354
rect 56802 119144 57554 119354
rect 57722 119144 58474 119354
rect 58642 119144 59394 119354
rect 59562 119144 60314 119354
rect 60482 119144 61234 119354
rect 61402 119144 62154 119354
rect 62322 119144 63074 119354
rect 63242 119144 63994 119354
rect 64162 119144 64914 119354
rect 65082 119144 65834 119354
rect 66002 119144 66754 119354
rect 66922 119144 67674 119354
rect 67842 119144 68594 119354
rect 68762 119144 69514 119354
rect 69682 119144 70434 119354
rect 70602 119144 71354 119354
rect 71522 119144 72274 119354
rect 72442 119144 73194 119354
rect 73362 119144 74114 119354
rect 74282 119144 75034 119354
rect 75202 119144 75954 119354
rect 76122 119144 76874 119354
rect 77042 119144 77794 119354
rect 77962 119144 78714 119354
rect 78882 119144 79634 119354
rect 79802 119144 80554 119354
rect 80722 119144 81474 119354
rect 81642 119144 82394 119354
rect 82562 119144 83314 119354
rect 83482 119144 84234 119354
rect 84402 119144 85154 119354
rect 85322 119144 86074 119354
rect 86242 119144 86994 119354
rect 87162 119144 87914 119354
rect 88082 119144 88834 119354
rect 89002 119144 89754 119354
rect 89922 119144 90674 119354
rect 90842 119144 91594 119354
rect 91762 119144 92514 119354
rect 92682 119144 93434 119354
rect 93602 119144 94354 119354
rect 94522 119144 95274 119354
rect 95442 119144 96194 119354
rect 96362 119144 97114 119354
rect 97282 119144 98034 119354
rect 98202 119144 98954 119354
rect 99122 119144 99874 119354
rect 100042 119144 100794 119354
rect 100962 119144 101714 119354
rect 101882 119144 102634 119354
rect 102802 119144 103554 119354
rect 103722 119144 104474 119354
rect 104642 119144 105394 119354
rect 105562 119144 106314 119354
rect 106482 119144 107234 119354
rect 107402 119144 108154 119354
rect 108322 119144 109074 119354
rect 109242 119144 109994 119354
rect 110162 119144 110914 119354
rect 111082 119144 111834 119354
rect 112002 119144 112754 119354
rect 112922 119144 113674 119354
rect 113842 119144 114594 119354
rect 114762 119144 115514 119354
rect 115682 119144 116434 119354
rect 116602 119144 117354 119354
rect 117522 119144 118274 119354
rect 118442 119144 119194 119354
rect 119362 119144 119764 119354
rect 480 856 119764 119144
rect 480 734 1434 856
rect 1602 734 2354 856
rect 2522 734 3274 856
rect 3442 734 4194 856
rect 4362 734 5114 856
rect 5282 734 6034 856
rect 6202 734 6954 856
rect 7122 734 7874 856
rect 8042 734 8794 856
rect 8962 734 9714 856
rect 9882 734 10634 856
rect 10802 734 11554 856
rect 11722 734 12474 856
rect 12642 734 13394 856
rect 13562 734 14314 856
rect 14482 734 15234 856
rect 15402 734 16154 856
rect 16322 734 17074 856
rect 17242 734 17994 856
rect 18162 734 18914 856
rect 19082 734 19834 856
rect 20002 734 20754 856
rect 20922 734 21674 856
rect 21842 734 22594 856
rect 22762 734 23514 856
rect 23682 734 24434 856
rect 24602 734 25354 856
rect 25522 734 26274 856
rect 26442 734 27194 856
rect 27362 734 28114 856
rect 28282 734 29034 856
rect 29202 734 29954 856
rect 30122 734 30874 856
rect 31042 734 31794 856
rect 31962 734 32714 856
rect 32882 734 33634 856
rect 33802 734 34554 856
rect 34722 734 35474 856
rect 35642 734 36394 856
rect 36562 734 37314 856
rect 37482 734 38234 856
rect 38402 734 39154 856
rect 39322 734 40074 856
rect 40242 734 40994 856
rect 41162 734 41914 856
rect 42082 734 42834 856
rect 43002 734 43754 856
rect 43922 734 44674 856
rect 44842 734 45594 856
rect 45762 734 46514 856
rect 46682 734 47434 856
rect 47602 734 48354 856
rect 48522 734 49274 856
rect 49442 734 50194 856
rect 50362 734 51114 856
rect 51282 734 52034 856
rect 52202 734 52954 856
rect 53122 734 53874 856
rect 54042 734 54794 856
rect 54962 734 55714 856
rect 55882 734 56634 856
rect 56802 734 57554 856
rect 57722 734 58474 856
rect 58642 734 59394 856
rect 59562 734 60314 856
rect 60482 734 61234 856
rect 61402 734 62154 856
rect 62322 734 63074 856
rect 63242 734 63994 856
rect 64162 734 64914 856
rect 65082 734 65834 856
rect 66002 734 66754 856
rect 66922 734 67674 856
rect 67842 734 68594 856
rect 68762 734 69514 856
rect 69682 734 70434 856
rect 70602 734 71354 856
rect 71522 734 72274 856
rect 72442 734 73194 856
rect 73362 734 74114 856
rect 74282 734 75034 856
rect 75202 734 75954 856
rect 76122 734 76874 856
rect 77042 734 77794 856
rect 77962 734 78714 856
rect 78882 734 79634 856
rect 79802 734 80554 856
rect 80722 734 81474 856
rect 81642 734 82394 856
rect 82562 734 83314 856
rect 83482 734 84234 856
rect 84402 734 85154 856
rect 85322 734 86074 856
rect 86242 734 86994 856
rect 87162 734 87914 856
rect 88082 734 88834 856
rect 89002 734 89754 856
rect 89922 734 90674 856
rect 90842 734 91594 856
rect 91762 734 92514 856
rect 92682 734 93434 856
rect 93602 734 94354 856
rect 94522 734 95274 856
rect 95442 734 96194 856
rect 96362 734 97114 856
rect 97282 734 98034 856
rect 98202 734 98954 856
rect 99122 734 99874 856
rect 100042 734 100794 856
rect 100962 734 101714 856
rect 101882 734 102634 856
rect 102802 734 103554 856
rect 103722 734 104474 856
rect 104642 734 105394 856
rect 105562 734 106314 856
rect 106482 734 107234 856
rect 107402 734 108154 856
rect 108322 734 109074 856
rect 109242 734 109994 856
rect 110162 734 110914 856
rect 111082 734 111834 856
rect 112002 734 112754 856
rect 112922 734 113674 856
rect 113842 734 114594 856
rect 114762 734 115514 856
rect 115682 734 116434 856
rect 116602 734 117354 856
rect 117522 734 118274 856
rect 118442 734 119764 856
<< metal3 >>
rect 119200 111664 120000 111784
rect 119200 110848 120000 110968
rect 119200 110032 120000 110152
rect 119200 109216 120000 109336
rect 119200 108400 120000 108520
rect 119200 107584 120000 107704
rect 119200 106768 120000 106888
rect 119200 105952 120000 106072
rect 119200 105136 120000 105256
rect 119200 104320 120000 104440
rect 119200 103504 120000 103624
rect 119200 102688 120000 102808
rect 119200 101872 120000 101992
rect 119200 101056 120000 101176
rect 119200 100240 120000 100360
rect 119200 99424 120000 99544
rect 119200 98608 120000 98728
rect 119200 97792 120000 97912
rect 119200 96976 120000 97096
rect 119200 96160 120000 96280
rect 119200 95344 120000 95464
rect 119200 94528 120000 94648
rect 119200 93712 120000 93832
rect 119200 92896 120000 93016
rect 119200 92080 120000 92200
rect 119200 91264 120000 91384
rect 119200 90448 120000 90568
rect 119200 89632 120000 89752
rect 119200 88816 120000 88936
rect 119200 88000 120000 88120
rect 119200 87184 120000 87304
rect 119200 86368 120000 86488
rect 119200 85552 120000 85672
rect 119200 84736 120000 84856
rect 119200 83920 120000 84040
rect 119200 83104 120000 83224
rect 119200 82288 120000 82408
rect 119200 81472 120000 81592
rect 119200 80656 120000 80776
rect 119200 79840 120000 79960
rect 119200 79024 120000 79144
rect 119200 78208 120000 78328
rect 119200 77392 120000 77512
rect 119200 76576 120000 76696
rect 119200 75760 120000 75880
rect 119200 74944 120000 75064
rect 119200 74128 120000 74248
rect 119200 73312 120000 73432
rect 119200 72496 120000 72616
rect 119200 71680 120000 71800
rect 119200 70864 120000 70984
rect 119200 70048 120000 70168
rect 119200 69232 120000 69352
rect 119200 68416 120000 68536
rect 119200 67600 120000 67720
rect 119200 66784 120000 66904
rect 119200 65968 120000 66088
rect 119200 65152 120000 65272
rect 119200 64336 120000 64456
rect 119200 63520 120000 63640
rect 119200 62704 120000 62824
rect 119200 61888 120000 62008
rect 119200 61072 120000 61192
rect 119200 60256 120000 60376
rect 119200 59440 120000 59560
rect 119200 58624 120000 58744
rect 119200 57808 120000 57928
rect 119200 56992 120000 57112
rect 119200 56176 120000 56296
rect 119200 55360 120000 55480
rect 119200 54544 120000 54664
rect 119200 53728 120000 53848
rect 119200 52912 120000 53032
rect 119200 52096 120000 52216
rect 119200 51280 120000 51400
rect 119200 50464 120000 50584
rect 119200 49648 120000 49768
rect 119200 48832 120000 48952
rect 119200 48016 120000 48136
rect 119200 47200 120000 47320
rect 119200 46384 120000 46504
rect 119200 45568 120000 45688
rect 119200 44752 120000 44872
rect 119200 43936 120000 44056
rect 119200 43120 120000 43240
rect 119200 42304 120000 42424
rect 119200 41488 120000 41608
rect 119200 40672 120000 40792
rect 119200 39856 120000 39976
rect 119200 39040 120000 39160
rect 119200 38224 120000 38344
rect 119200 37408 120000 37528
rect 119200 36592 120000 36712
rect 119200 35776 120000 35896
rect 119200 34960 120000 35080
rect 119200 34144 120000 34264
rect 119200 33328 120000 33448
rect 119200 32512 120000 32632
rect 119200 31696 120000 31816
rect 119200 30880 120000 31000
rect 119200 30064 120000 30184
rect 119200 29248 120000 29368
rect 119200 28432 120000 28552
rect 119200 27616 120000 27736
rect 119200 26800 120000 26920
rect 119200 25984 120000 26104
rect 119200 25168 120000 25288
rect 119200 24352 120000 24472
rect 119200 23536 120000 23656
rect 119200 22720 120000 22840
rect 119200 21904 120000 22024
rect 119200 21088 120000 21208
rect 119200 20272 120000 20392
rect 119200 19456 120000 19576
rect 119200 18640 120000 18760
rect 119200 17824 120000 17944
rect 119200 17008 120000 17128
rect 119200 16192 120000 16312
rect 119200 15376 120000 15496
rect 119200 14560 120000 14680
rect 119200 13744 120000 13864
rect 119200 12928 120000 13048
rect 119200 12112 120000 12232
rect 119200 11296 120000 11416
rect 119200 10480 120000 10600
rect 119200 9664 120000 9784
rect 119200 8848 120000 8968
rect 119200 8032 120000 8152
<< obsm3 >>
rect 657 111864 119495 117537
rect 657 111584 119120 111864
rect 657 111048 119495 111584
rect 657 110768 119120 111048
rect 657 110232 119495 110768
rect 657 109952 119120 110232
rect 657 109416 119495 109952
rect 657 109136 119120 109416
rect 657 108600 119495 109136
rect 657 108320 119120 108600
rect 657 107784 119495 108320
rect 657 107504 119120 107784
rect 657 106968 119495 107504
rect 657 106688 119120 106968
rect 657 106152 119495 106688
rect 657 105872 119120 106152
rect 657 105336 119495 105872
rect 657 105056 119120 105336
rect 657 104520 119495 105056
rect 657 104240 119120 104520
rect 657 103704 119495 104240
rect 657 103424 119120 103704
rect 657 102888 119495 103424
rect 657 102608 119120 102888
rect 657 102072 119495 102608
rect 657 101792 119120 102072
rect 657 101256 119495 101792
rect 657 100976 119120 101256
rect 657 100440 119495 100976
rect 657 100160 119120 100440
rect 657 99624 119495 100160
rect 657 99344 119120 99624
rect 657 98808 119495 99344
rect 657 98528 119120 98808
rect 657 97992 119495 98528
rect 657 97712 119120 97992
rect 657 97176 119495 97712
rect 657 96896 119120 97176
rect 657 96360 119495 96896
rect 657 96080 119120 96360
rect 657 95544 119495 96080
rect 657 95264 119120 95544
rect 657 94728 119495 95264
rect 657 94448 119120 94728
rect 657 93912 119495 94448
rect 657 93632 119120 93912
rect 657 93096 119495 93632
rect 657 92816 119120 93096
rect 657 92280 119495 92816
rect 657 92000 119120 92280
rect 657 91464 119495 92000
rect 657 91184 119120 91464
rect 657 90648 119495 91184
rect 657 90368 119120 90648
rect 657 89832 119495 90368
rect 657 89552 119120 89832
rect 657 89016 119495 89552
rect 657 88736 119120 89016
rect 657 88200 119495 88736
rect 657 87920 119120 88200
rect 657 87384 119495 87920
rect 657 87104 119120 87384
rect 657 86568 119495 87104
rect 657 86288 119120 86568
rect 657 85752 119495 86288
rect 657 85472 119120 85752
rect 657 84936 119495 85472
rect 657 84656 119120 84936
rect 657 84120 119495 84656
rect 657 83840 119120 84120
rect 657 83304 119495 83840
rect 657 83024 119120 83304
rect 657 82488 119495 83024
rect 657 82208 119120 82488
rect 657 81672 119495 82208
rect 657 81392 119120 81672
rect 657 80856 119495 81392
rect 657 80576 119120 80856
rect 657 80040 119495 80576
rect 657 79760 119120 80040
rect 657 79224 119495 79760
rect 657 78944 119120 79224
rect 657 78408 119495 78944
rect 657 78128 119120 78408
rect 657 77592 119495 78128
rect 657 77312 119120 77592
rect 657 76776 119495 77312
rect 657 76496 119120 76776
rect 657 75960 119495 76496
rect 657 75680 119120 75960
rect 657 75144 119495 75680
rect 657 74864 119120 75144
rect 657 74328 119495 74864
rect 657 74048 119120 74328
rect 657 73512 119495 74048
rect 657 73232 119120 73512
rect 657 72696 119495 73232
rect 657 72416 119120 72696
rect 657 71880 119495 72416
rect 657 71600 119120 71880
rect 657 71064 119495 71600
rect 657 70784 119120 71064
rect 657 70248 119495 70784
rect 657 69968 119120 70248
rect 657 69432 119495 69968
rect 657 69152 119120 69432
rect 657 68616 119495 69152
rect 657 68336 119120 68616
rect 657 67800 119495 68336
rect 657 67520 119120 67800
rect 657 66984 119495 67520
rect 657 66704 119120 66984
rect 657 66168 119495 66704
rect 657 65888 119120 66168
rect 657 65352 119495 65888
rect 657 65072 119120 65352
rect 657 64536 119495 65072
rect 657 64256 119120 64536
rect 657 63720 119495 64256
rect 657 63440 119120 63720
rect 657 62904 119495 63440
rect 657 62624 119120 62904
rect 657 62088 119495 62624
rect 657 61808 119120 62088
rect 657 61272 119495 61808
rect 657 60992 119120 61272
rect 657 60456 119495 60992
rect 657 60176 119120 60456
rect 657 59640 119495 60176
rect 657 59360 119120 59640
rect 657 58824 119495 59360
rect 657 58544 119120 58824
rect 657 58008 119495 58544
rect 657 57728 119120 58008
rect 657 57192 119495 57728
rect 657 56912 119120 57192
rect 657 56376 119495 56912
rect 657 56096 119120 56376
rect 657 55560 119495 56096
rect 657 55280 119120 55560
rect 657 54744 119495 55280
rect 657 54464 119120 54744
rect 657 53928 119495 54464
rect 657 53648 119120 53928
rect 657 53112 119495 53648
rect 657 52832 119120 53112
rect 657 52296 119495 52832
rect 657 52016 119120 52296
rect 657 51480 119495 52016
rect 657 51200 119120 51480
rect 657 50664 119495 51200
rect 657 50384 119120 50664
rect 657 49848 119495 50384
rect 657 49568 119120 49848
rect 657 49032 119495 49568
rect 657 48752 119120 49032
rect 657 48216 119495 48752
rect 657 47936 119120 48216
rect 657 47400 119495 47936
rect 657 47120 119120 47400
rect 657 46584 119495 47120
rect 657 46304 119120 46584
rect 657 45768 119495 46304
rect 657 45488 119120 45768
rect 657 44952 119495 45488
rect 657 44672 119120 44952
rect 657 44136 119495 44672
rect 657 43856 119120 44136
rect 657 43320 119495 43856
rect 657 43040 119120 43320
rect 657 42504 119495 43040
rect 657 42224 119120 42504
rect 657 41688 119495 42224
rect 657 41408 119120 41688
rect 657 40872 119495 41408
rect 657 40592 119120 40872
rect 657 40056 119495 40592
rect 657 39776 119120 40056
rect 657 39240 119495 39776
rect 657 38960 119120 39240
rect 657 38424 119495 38960
rect 657 38144 119120 38424
rect 657 37608 119495 38144
rect 657 37328 119120 37608
rect 657 36792 119495 37328
rect 657 36512 119120 36792
rect 657 35976 119495 36512
rect 657 35696 119120 35976
rect 657 35160 119495 35696
rect 657 34880 119120 35160
rect 657 34344 119495 34880
rect 657 34064 119120 34344
rect 657 33528 119495 34064
rect 657 33248 119120 33528
rect 657 32712 119495 33248
rect 657 32432 119120 32712
rect 657 31896 119495 32432
rect 657 31616 119120 31896
rect 657 31080 119495 31616
rect 657 30800 119120 31080
rect 657 30264 119495 30800
rect 657 29984 119120 30264
rect 657 29448 119495 29984
rect 657 29168 119120 29448
rect 657 28632 119495 29168
rect 657 28352 119120 28632
rect 657 27816 119495 28352
rect 657 27536 119120 27816
rect 657 27000 119495 27536
rect 657 26720 119120 27000
rect 657 26184 119495 26720
rect 657 25904 119120 26184
rect 657 25368 119495 25904
rect 657 25088 119120 25368
rect 657 24552 119495 25088
rect 657 24272 119120 24552
rect 657 23736 119495 24272
rect 657 23456 119120 23736
rect 657 22920 119495 23456
rect 657 22640 119120 22920
rect 657 22104 119495 22640
rect 657 21824 119120 22104
rect 657 21288 119495 21824
rect 657 21008 119120 21288
rect 657 20472 119495 21008
rect 657 20192 119120 20472
rect 657 19656 119495 20192
rect 657 19376 119120 19656
rect 657 18840 119495 19376
rect 657 18560 119120 18840
rect 657 18024 119495 18560
rect 657 17744 119120 18024
rect 657 17208 119495 17744
rect 657 16928 119120 17208
rect 657 16392 119495 16928
rect 657 16112 119120 16392
rect 657 15576 119495 16112
rect 657 15296 119120 15576
rect 657 14760 119495 15296
rect 657 14480 119120 14760
rect 657 13944 119495 14480
rect 657 13664 119120 13944
rect 657 13128 119495 13664
rect 657 12848 119120 13128
rect 657 12312 119495 12848
rect 657 12032 119120 12312
rect 657 11496 119495 12032
rect 657 11216 119120 11496
rect 657 10680 119495 11216
rect 657 10400 119120 10680
rect 657 9864 119495 10400
rect 657 9584 119120 9864
rect 657 9048 119495 9584
rect 657 8768 119120 9048
rect 657 8232 119495 8768
rect 657 7952 119120 8232
rect 657 1803 119495 7952
<< metal4 >>
rect 1794 2128 2414 117552
rect 19794 2128 20414 117552
rect 37794 2128 38414 117552
rect 55794 2128 56414 117552
rect 73794 2128 74414 117552
rect 91794 2128 92414 117552
rect 109794 2128 110414 117552
<< obsm4 >>
rect 1531 2048 1714 112029
rect 2494 2048 19714 112029
rect 20494 2048 37714 112029
rect 38494 2048 55714 112029
rect 56494 2048 73714 112029
rect 74494 2048 91714 112029
rect 92494 2048 109714 112029
rect 110494 2048 116781 112029
rect 1531 1803 116781 2048
<< labels >>
rlabel metal4 s 19794 2128 20414 117552 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 55794 2128 56414 117552 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 91794 2128 92414 117552 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1794 2128 2414 117552 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 37794 2128 38414 117552 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 73794 2128 74414 117552 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 109794 2128 110414 117552 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 119200 8032 120000 8152 6 a[0]
port 3 nsew signal input
rlabel metal3 s 119200 16192 120000 16312 6 a[10]
port 4 nsew signal input
rlabel metal3 s 119200 17008 120000 17128 6 a[11]
port 5 nsew signal input
rlabel metal3 s 119200 17824 120000 17944 6 a[12]
port 6 nsew signal input
rlabel metal3 s 119200 18640 120000 18760 6 a[13]
port 7 nsew signal input
rlabel metal3 s 119200 19456 120000 19576 6 a[14]
port 8 nsew signal input
rlabel metal3 s 119200 20272 120000 20392 6 a[15]
port 9 nsew signal input
rlabel metal3 s 119200 21088 120000 21208 6 a[16]
port 10 nsew signal input
rlabel metal3 s 119200 21904 120000 22024 6 a[17]
port 11 nsew signal input
rlabel metal3 s 119200 22720 120000 22840 6 a[18]
port 12 nsew signal input
rlabel metal3 s 119200 23536 120000 23656 6 a[19]
port 13 nsew signal input
rlabel metal3 s 119200 8848 120000 8968 6 a[1]
port 14 nsew signal input
rlabel metal3 s 119200 24352 120000 24472 6 a[20]
port 15 nsew signal input
rlabel metal3 s 119200 25168 120000 25288 6 a[21]
port 16 nsew signal input
rlabel metal3 s 119200 25984 120000 26104 6 a[22]
port 17 nsew signal input
rlabel metal3 s 119200 26800 120000 26920 6 a[23]
port 18 nsew signal input
rlabel metal3 s 119200 27616 120000 27736 6 a[24]
port 19 nsew signal input
rlabel metal3 s 119200 28432 120000 28552 6 a[25]
port 20 nsew signal input
rlabel metal3 s 119200 29248 120000 29368 6 a[26]
port 21 nsew signal input
rlabel metal3 s 119200 30064 120000 30184 6 a[27]
port 22 nsew signal input
rlabel metal3 s 119200 30880 120000 31000 6 a[28]
port 23 nsew signal input
rlabel metal3 s 119200 31696 120000 31816 6 a[29]
port 24 nsew signal input
rlabel metal3 s 119200 9664 120000 9784 6 a[2]
port 25 nsew signal input
rlabel metal3 s 119200 32512 120000 32632 6 a[30]
port 26 nsew signal input
rlabel metal3 s 119200 33328 120000 33448 6 a[31]
port 27 nsew signal input
rlabel metal3 s 119200 34144 120000 34264 6 a[32]
port 28 nsew signal input
rlabel metal3 s 119200 34960 120000 35080 6 a[33]
port 29 nsew signal input
rlabel metal3 s 119200 35776 120000 35896 6 a[34]
port 30 nsew signal input
rlabel metal3 s 119200 36592 120000 36712 6 a[35]
port 31 nsew signal input
rlabel metal3 s 119200 37408 120000 37528 6 a[36]
port 32 nsew signal input
rlabel metal3 s 119200 38224 120000 38344 6 a[37]
port 33 nsew signal input
rlabel metal3 s 119200 39040 120000 39160 6 a[38]
port 34 nsew signal input
rlabel metal3 s 119200 39856 120000 39976 6 a[39]
port 35 nsew signal input
rlabel metal3 s 119200 10480 120000 10600 6 a[3]
port 36 nsew signal input
rlabel metal3 s 119200 40672 120000 40792 6 a[40]
port 37 nsew signal input
rlabel metal3 s 119200 41488 120000 41608 6 a[41]
port 38 nsew signal input
rlabel metal3 s 119200 42304 120000 42424 6 a[42]
port 39 nsew signal input
rlabel metal3 s 119200 43120 120000 43240 6 a[43]
port 40 nsew signal input
rlabel metal3 s 119200 43936 120000 44056 6 a[44]
port 41 nsew signal input
rlabel metal3 s 119200 44752 120000 44872 6 a[45]
port 42 nsew signal input
rlabel metal3 s 119200 45568 120000 45688 6 a[46]
port 43 nsew signal input
rlabel metal3 s 119200 46384 120000 46504 6 a[47]
port 44 nsew signal input
rlabel metal3 s 119200 47200 120000 47320 6 a[48]
port 45 nsew signal input
rlabel metal3 s 119200 48016 120000 48136 6 a[49]
port 46 nsew signal input
rlabel metal3 s 119200 11296 120000 11416 6 a[4]
port 47 nsew signal input
rlabel metal3 s 119200 48832 120000 48952 6 a[50]
port 48 nsew signal input
rlabel metal3 s 119200 49648 120000 49768 6 a[51]
port 49 nsew signal input
rlabel metal3 s 119200 50464 120000 50584 6 a[52]
port 50 nsew signal input
rlabel metal3 s 119200 51280 120000 51400 6 a[53]
port 51 nsew signal input
rlabel metal3 s 119200 52096 120000 52216 6 a[54]
port 52 nsew signal input
rlabel metal3 s 119200 52912 120000 53032 6 a[55]
port 53 nsew signal input
rlabel metal3 s 119200 53728 120000 53848 6 a[56]
port 54 nsew signal input
rlabel metal3 s 119200 54544 120000 54664 6 a[57]
port 55 nsew signal input
rlabel metal3 s 119200 55360 120000 55480 6 a[58]
port 56 nsew signal input
rlabel metal3 s 119200 56176 120000 56296 6 a[59]
port 57 nsew signal input
rlabel metal3 s 119200 12112 120000 12232 6 a[5]
port 58 nsew signal input
rlabel metal3 s 119200 56992 120000 57112 6 a[60]
port 59 nsew signal input
rlabel metal3 s 119200 57808 120000 57928 6 a[61]
port 60 nsew signal input
rlabel metal3 s 119200 58624 120000 58744 6 a[62]
port 61 nsew signal input
rlabel metal3 s 119200 59440 120000 59560 6 a[63]
port 62 nsew signal input
rlabel metal3 s 119200 12928 120000 13048 6 a[6]
port 63 nsew signal input
rlabel metal3 s 119200 13744 120000 13864 6 a[7]
port 64 nsew signal input
rlabel metal3 s 119200 14560 120000 14680 6 a[8]
port 65 nsew signal input
rlabel metal3 s 119200 15376 120000 15496 6 a[9]
port 66 nsew signal input
rlabel metal3 s 119200 60256 120000 60376 6 b[0]
port 67 nsew signal input
rlabel metal3 s 119200 68416 120000 68536 6 b[10]
port 68 nsew signal input
rlabel metal3 s 119200 69232 120000 69352 6 b[11]
port 69 nsew signal input
rlabel metal3 s 119200 70048 120000 70168 6 b[12]
port 70 nsew signal input
rlabel metal3 s 119200 70864 120000 70984 6 b[13]
port 71 nsew signal input
rlabel metal3 s 119200 71680 120000 71800 6 b[14]
port 72 nsew signal input
rlabel metal3 s 119200 72496 120000 72616 6 b[15]
port 73 nsew signal input
rlabel metal3 s 119200 73312 120000 73432 6 b[16]
port 74 nsew signal input
rlabel metal3 s 119200 74128 120000 74248 6 b[17]
port 75 nsew signal input
rlabel metal3 s 119200 74944 120000 75064 6 b[18]
port 76 nsew signal input
rlabel metal3 s 119200 75760 120000 75880 6 b[19]
port 77 nsew signal input
rlabel metal3 s 119200 61072 120000 61192 6 b[1]
port 78 nsew signal input
rlabel metal3 s 119200 76576 120000 76696 6 b[20]
port 79 nsew signal input
rlabel metal3 s 119200 77392 120000 77512 6 b[21]
port 80 nsew signal input
rlabel metal3 s 119200 78208 120000 78328 6 b[22]
port 81 nsew signal input
rlabel metal3 s 119200 79024 120000 79144 6 b[23]
port 82 nsew signal input
rlabel metal3 s 119200 79840 120000 79960 6 b[24]
port 83 nsew signal input
rlabel metal3 s 119200 80656 120000 80776 6 b[25]
port 84 nsew signal input
rlabel metal3 s 119200 81472 120000 81592 6 b[26]
port 85 nsew signal input
rlabel metal3 s 119200 82288 120000 82408 6 b[27]
port 86 nsew signal input
rlabel metal3 s 119200 83104 120000 83224 6 b[28]
port 87 nsew signal input
rlabel metal3 s 119200 83920 120000 84040 6 b[29]
port 88 nsew signal input
rlabel metal3 s 119200 61888 120000 62008 6 b[2]
port 89 nsew signal input
rlabel metal3 s 119200 84736 120000 84856 6 b[30]
port 90 nsew signal input
rlabel metal3 s 119200 85552 120000 85672 6 b[31]
port 91 nsew signal input
rlabel metal3 s 119200 86368 120000 86488 6 b[32]
port 92 nsew signal input
rlabel metal3 s 119200 87184 120000 87304 6 b[33]
port 93 nsew signal input
rlabel metal3 s 119200 88000 120000 88120 6 b[34]
port 94 nsew signal input
rlabel metal3 s 119200 88816 120000 88936 6 b[35]
port 95 nsew signal input
rlabel metal3 s 119200 89632 120000 89752 6 b[36]
port 96 nsew signal input
rlabel metal3 s 119200 90448 120000 90568 6 b[37]
port 97 nsew signal input
rlabel metal3 s 119200 91264 120000 91384 6 b[38]
port 98 nsew signal input
rlabel metal3 s 119200 92080 120000 92200 6 b[39]
port 99 nsew signal input
rlabel metal3 s 119200 62704 120000 62824 6 b[3]
port 100 nsew signal input
rlabel metal3 s 119200 92896 120000 93016 6 b[40]
port 101 nsew signal input
rlabel metal3 s 119200 93712 120000 93832 6 b[41]
port 102 nsew signal input
rlabel metal3 s 119200 94528 120000 94648 6 b[42]
port 103 nsew signal input
rlabel metal3 s 119200 95344 120000 95464 6 b[43]
port 104 nsew signal input
rlabel metal3 s 119200 96160 120000 96280 6 b[44]
port 105 nsew signal input
rlabel metal3 s 119200 96976 120000 97096 6 b[45]
port 106 nsew signal input
rlabel metal3 s 119200 97792 120000 97912 6 b[46]
port 107 nsew signal input
rlabel metal3 s 119200 98608 120000 98728 6 b[47]
port 108 nsew signal input
rlabel metal3 s 119200 99424 120000 99544 6 b[48]
port 109 nsew signal input
rlabel metal3 s 119200 100240 120000 100360 6 b[49]
port 110 nsew signal input
rlabel metal3 s 119200 63520 120000 63640 6 b[4]
port 111 nsew signal input
rlabel metal3 s 119200 101056 120000 101176 6 b[50]
port 112 nsew signal input
rlabel metal3 s 119200 101872 120000 101992 6 b[51]
port 113 nsew signal input
rlabel metal3 s 119200 102688 120000 102808 6 b[52]
port 114 nsew signal input
rlabel metal3 s 119200 103504 120000 103624 6 b[53]
port 115 nsew signal input
rlabel metal3 s 119200 104320 120000 104440 6 b[54]
port 116 nsew signal input
rlabel metal3 s 119200 105136 120000 105256 6 b[55]
port 117 nsew signal input
rlabel metal3 s 119200 105952 120000 106072 6 b[56]
port 118 nsew signal input
rlabel metal3 s 119200 106768 120000 106888 6 b[57]
port 119 nsew signal input
rlabel metal3 s 119200 107584 120000 107704 6 b[58]
port 120 nsew signal input
rlabel metal3 s 119200 108400 120000 108520 6 b[59]
port 121 nsew signal input
rlabel metal3 s 119200 64336 120000 64456 6 b[5]
port 122 nsew signal input
rlabel metal3 s 119200 109216 120000 109336 6 b[60]
port 123 nsew signal input
rlabel metal3 s 119200 110032 120000 110152 6 b[61]
port 124 nsew signal input
rlabel metal3 s 119200 110848 120000 110968 6 b[62]
port 125 nsew signal input
rlabel metal3 s 119200 111664 120000 111784 6 b[63]
port 126 nsew signal input
rlabel metal3 s 119200 65152 120000 65272 6 b[6]
port 127 nsew signal input
rlabel metal3 s 119200 65968 120000 66088 6 b[7]
port 128 nsew signal input
rlabel metal3 s 119200 66784 120000 66904 6 b[8]
port 129 nsew signal input
rlabel metal3 s 119200 67600 120000 67720 6 b[9]
port 130 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 c[0]
port 131 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 c[100]
port 132 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 c[101]
port 133 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 c[102]
port 134 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 c[103]
port 135 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 c[104]
port 136 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 c[105]
port 137 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 c[106]
port 138 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 c[107]
port 139 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 c[108]
port 140 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 c[109]
port 141 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 c[10]
port 142 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 c[110]
port 143 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 c[111]
port 144 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 c[112]
port 145 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 c[113]
port 146 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 c[114]
port 147 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 c[115]
port 148 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 c[116]
port 149 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 c[117]
port 150 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 c[118]
port 151 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 c[119]
port 152 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 c[11]
port 153 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 c[120]
port 154 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 c[121]
port 155 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 c[122]
port 156 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 c[123]
port 157 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 c[124]
port 158 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 c[125]
port 159 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 c[126]
port 160 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 c[127]
port 161 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 c[12]
port 162 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 c[13]
port 163 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 c[14]
port 164 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 c[15]
port 165 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 c[16]
port 166 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 c[17]
port 167 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 c[18]
port 168 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 c[19]
port 169 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 c[1]
port 170 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 c[20]
port 171 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 c[21]
port 172 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 c[22]
port 173 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 c[23]
port 174 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 c[24]
port 175 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 c[25]
port 176 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 c[26]
port 177 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 c[27]
port 178 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 c[28]
port 179 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 c[29]
port 180 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 c[2]
port 181 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 c[30]
port 182 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 c[31]
port 183 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 c[32]
port 184 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 c[33]
port 185 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 c[34]
port 186 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 c[35]
port 187 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 c[36]
port 188 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 c[37]
port 189 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 c[38]
port 190 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 c[39]
port 191 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 c[3]
port 192 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 c[40]
port 193 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 c[41]
port 194 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 c[42]
port 195 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 c[43]
port 196 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 c[44]
port 197 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 c[45]
port 198 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 c[46]
port 199 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 c[47]
port 200 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 c[48]
port 201 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 c[49]
port 202 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 c[4]
port 203 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 c[50]
port 204 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 c[51]
port 205 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 c[52]
port 206 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 c[53]
port 207 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 c[54]
port 208 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 c[55]
port 209 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 c[56]
port 210 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 c[57]
port 211 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 c[58]
port 212 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 c[59]
port 213 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 c[5]
port 214 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 c[60]
port 215 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 c[61]
port 216 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 c[62]
port 217 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 c[63]
port 218 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 c[64]
port 219 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 c[65]
port 220 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 c[66]
port 221 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 c[67]
port 222 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 c[68]
port 223 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 c[69]
port 224 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 c[6]
port 225 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 c[70]
port 226 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 c[71]
port 227 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 c[72]
port 228 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 c[73]
port 229 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 c[74]
port 230 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 c[75]
port 231 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 c[76]
port 232 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 c[77]
port 233 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 c[78]
port 234 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 c[79]
port 235 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 c[7]
port 236 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 c[80]
port 237 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 c[81]
port 238 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 c[82]
port 239 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 c[83]
port 240 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 c[84]
port 241 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 c[85]
port 242 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 c[86]
port 243 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 c[87]
port 244 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 c[88]
port 245 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 c[89]
port 246 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 c[8]
port 247 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 c[90]
port 248 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 c[91]
port 249 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 c[92]
port 250 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 c[93]
port 251 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 c[94]
port 252 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 c[95]
port 253 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 c[96]
port 254 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 c[97]
port 255 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 c[98]
port 256 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 c[99]
port 257 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 c[9]
port 258 nsew signal input
rlabel metal2 s 119250 119200 119306 120000 6 clk
port 259 nsew signal input
rlabel metal2 s 570 119200 626 120000 6 o[0]
port 260 nsew signal output
rlabel metal2 s 92570 119200 92626 120000 6 o[100]
port 261 nsew signal output
rlabel metal2 s 93490 119200 93546 120000 6 o[101]
port 262 nsew signal output
rlabel metal2 s 94410 119200 94466 120000 6 o[102]
port 263 nsew signal output
rlabel metal2 s 95330 119200 95386 120000 6 o[103]
port 264 nsew signal output
rlabel metal2 s 96250 119200 96306 120000 6 o[104]
port 265 nsew signal output
rlabel metal2 s 97170 119200 97226 120000 6 o[105]
port 266 nsew signal output
rlabel metal2 s 98090 119200 98146 120000 6 o[106]
port 267 nsew signal output
rlabel metal2 s 99010 119200 99066 120000 6 o[107]
port 268 nsew signal output
rlabel metal2 s 99930 119200 99986 120000 6 o[108]
port 269 nsew signal output
rlabel metal2 s 100850 119200 100906 120000 6 o[109]
port 270 nsew signal output
rlabel metal2 s 9770 119200 9826 120000 6 o[10]
port 271 nsew signal output
rlabel metal2 s 101770 119200 101826 120000 6 o[110]
port 272 nsew signal output
rlabel metal2 s 102690 119200 102746 120000 6 o[111]
port 273 nsew signal output
rlabel metal2 s 103610 119200 103666 120000 6 o[112]
port 274 nsew signal output
rlabel metal2 s 104530 119200 104586 120000 6 o[113]
port 275 nsew signal output
rlabel metal2 s 105450 119200 105506 120000 6 o[114]
port 276 nsew signal output
rlabel metal2 s 106370 119200 106426 120000 6 o[115]
port 277 nsew signal output
rlabel metal2 s 107290 119200 107346 120000 6 o[116]
port 278 nsew signal output
rlabel metal2 s 108210 119200 108266 120000 6 o[117]
port 279 nsew signal output
rlabel metal2 s 109130 119200 109186 120000 6 o[118]
port 280 nsew signal output
rlabel metal2 s 110050 119200 110106 120000 6 o[119]
port 281 nsew signal output
rlabel metal2 s 10690 119200 10746 120000 6 o[11]
port 282 nsew signal output
rlabel metal2 s 110970 119200 111026 120000 6 o[120]
port 283 nsew signal output
rlabel metal2 s 111890 119200 111946 120000 6 o[121]
port 284 nsew signal output
rlabel metal2 s 112810 119200 112866 120000 6 o[122]
port 285 nsew signal output
rlabel metal2 s 113730 119200 113786 120000 6 o[123]
port 286 nsew signal output
rlabel metal2 s 114650 119200 114706 120000 6 o[124]
port 287 nsew signal output
rlabel metal2 s 115570 119200 115626 120000 6 o[125]
port 288 nsew signal output
rlabel metal2 s 116490 119200 116546 120000 6 o[126]
port 289 nsew signal output
rlabel metal2 s 117410 119200 117466 120000 6 o[127]
port 290 nsew signal output
rlabel metal2 s 11610 119200 11666 120000 6 o[12]
port 291 nsew signal output
rlabel metal2 s 12530 119200 12586 120000 6 o[13]
port 292 nsew signal output
rlabel metal2 s 13450 119200 13506 120000 6 o[14]
port 293 nsew signal output
rlabel metal2 s 14370 119200 14426 120000 6 o[15]
port 294 nsew signal output
rlabel metal2 s 15290 119200 15346 120000 6 o[16]
port 295 nsew signal output
rlabel metal2 s 16210 119200 16266 120000 6 o[17]
port 296 nsew signal output
rlabel metal2 s 17130 119200 17186 120000 6 o[18]
port 297 nsew signal output
rlabel metal2 s 18050 119200 18106 120000 6 o[19]
port 298 nsew signal output
rlabel metal2 s 1490 119200 1546 120000 6 o[1]
port 299 nsew signal output
rlabel metal2 s 18970 119200 19026 120000 6 o[20]
port 300 nsew signal output
rlabel metal2 s 19890 119200 19946 120000 6 o[21]
port 301 nsew signal output
rlabel metal2 s 20810 119200 20866 120000 6 o[22]
port 302 nsew signal output
rlabel metal2 s 21730 119200 21786 120000 6 o[23]
port 303 nsew signal output
rlabel metal2 s 22650 119200 22706 120000 6 o[24]
port 304 nsew signal output
rlabel metal2 s 23570 119200 23626 120000 6 o[25]
port 305 nsew signal output
rlabel metal2 s 24490 119200 24546 120000 6 o[26]
port 306 nsew signal output
rlabel metal2 s 25410 119200 25466 120000 6 o[27]
port 307 nsew signal output
rlabel metal2 s 26330 119200 26386 120000 6 o[28]
port 308 nsew signal output
rlabel metal2 s 27250 119200 27306 120000 6 o[29]
port 309 nsew signal output
rlabel metal2 s 2410 119200 2466 120000 6 o[2]
port 310 nsew signal output
rlabel metal2 s 28170 119200 28226 120000 6 o[30]
port 311 nsew signal output
rlabel metal2 s 29090 119200 29146 120000 6 o[31]
port 312 nsew signal output
rlabel metal2 s 30010 119200 30066 120000 6 o[32]
port 313 nsew signal output
rlabel metal2 s 30930 119200 30986 120000 6 o[33]
port 314 nsew signal output
rlabel metal2 s 31850 119200 31906 120000 6 o[34]
port 315 nsew signal output
rlabel metal2 s 32770 119200 32826 120000 6 o[35]
port 316 nsew signal output
rlabel metal2 s 33690 119200 33746 120000 6 o[36]
port 317 nsew signal output
rlabel metal2 s 34610 119200 34666 120000 6 o[37]
port 318 nsew signal output
rlabel metal2 s 35530 119200 35586 120000 6 o[38]
port 319 nsew signal output
rlabel metal2 s 36450 119200 36506 120000 6 o[39]
port 320 nsew signal output
rlabel metal2 s 3330 119200 3386 120000 6 o[3]
port 321 nsew signal output
rlabel metal2 s 37370 119200 37426 120000 6 o[40]
port 322 nsew signal output
rlabel metal2 s 38290 119200 38346 120000 6 o[41]
port 323 nsew signal output
rlabel metal2 s 39210 119200 39266 120000 6 o[42]
port 324 nsew signal output
rlabel metal2 s 40130 119200 40186 120000 6 o[43]
port 325 nsew signal output
rlabel metal2 s 41050 119200 41106 120000 6 o[44]
port 326 nsew signal output
rlabel metal2 s 41970 119200 42026 120000 6 o[45]
port 327 nsew signal output
rlabel metal2 s 42890 119200 42946 120000 6 o[46]
port 328 nsew signal output
rlabel metal2 s 43810 119200 43866 120000 6 o[47]
port 329 nsew signal output
rlabel metal2 s 44730 119200 44786 120000 6 o[48]
port 330 nsew signal output
rlabel metal2 s 45650 119200 45706 120000 6 o[49]
port 331 nsew signal output
rlabel metal2 s 4250 119200 4306 120000 6 o[4]
port 332 nsew signal output
rlabel metal2 s 46570 119200 46626 120000 6 o[50]
port 333 nsew signal output
rlabel metal2 s 47490 119200 47546 120000 6 o[51]
port 334 nsew signal output
rlabel metal2 s 48410 119200 48466 120000 6 o[52]
port 335 nsew signal output
rlabel metal2 s 49330 119200 49386 120000 6 o[53]
port 336 nsew signal output
rlabel metal2 s 50250 119200 50306 120000 6 o[54]
port 337 nsew signal output
rlabel metal2 s 51170 119200 51226 120000 6 o[55]
port 338 nsew signal output
rlabel metal2 s 52090 119200 52146 120000 6 o[56]
port 339 nsew signal output
rlabel metal2 s 53010 119200 53066 120000 6 o[57]
port 340 nsew signal output
rlabel metal2 s 53930 119200 53986 120000 6 o[58]
port 341 nsew signal output
rlabel metal2 s 54850 119200 54906 120000 6 o[59]
port 342 nsew signal output
rlabel metal2 s 5170 119200 5226 120000 6 o[5]
port 343 nsew signal output
rlabel metal2 s 55770 119200 55826 120000 6 o[60]
port 344 nsew signal output
rlabel metal2 s 56690 119200 56746 120000 6 o[61]
port 345 nsew signal output
rlabel metal2 s 57610 119200 57666 120000 6 o[62]
port 346 nsew signal output
rlabel metal2 s 58530 119200 58586 120000 6 o[63]
port 347 nsew signal output
rlabel metal2 s 59450 119200 59506 120000 6 o[64]
port 348 nsew signal output
rlabel metal2 s 60370 119200 60426 120000 6 o[65]
port 349 nsew signal output
rlabel metal2 s 61290 119200 61346 120000 6 o[66]
port 350 nsew signal output
rlabel metal2 s 62210 119200 62266 120000 6 o[67]
port 351 nsew signal output
rlabel metal2 s 63130 119200 63186 120000 6 o[68]
port 352 nsew signal output
rlabel metal2 s 64050 119200 64106 120000 6 o[69]
port 353 nsew signal output
rlabel metal2 s 6090 119200 6146 120000 6 o[6]
port 354 nsew signal output
rlabel metal2 s 64970 119200 65026 120000 6 o[70]
port 355 nsew signal output
rlabel metal2 s 65890 119200 65946 120000 6 o[71]
port 356 nsew signal output
rlabel metal2 s 66810 119200 66866 120000 6 o[72]
port 357 nsew signal output
rlabel metal2 s 67730 119200 67786 120000 6 o[73]
port 358 nsew signal output
rlabel metal2 s 68650 119200 68706 120000 6 o[74]
port 359 nsew signal output
rlabel metal2 s 69570 119200 69626 120000 6 o[75]
port 360 nsew signal output
rlabel metal2 s 70490 119200 70546 120000 6 o[76]
port 361 nsew signal output
rlabel metal2 s 71410 119200 71466 120000 6 o[77]
port 362 nsew signal output
rlabel metal2 s 72330 119200 72386 120000 6 o[78]
port 363 nsew signal output
rlabel metal2 s 73250 119200 73306 120000 6 o[79]
port 364 nsew signal output
rlabel metal2 s 7010 119200 7066 120000 6 o[7]
port 365 nsew signal output
rlabel metal2 s 74170 119200 74226 120000 6 o[80]
port 366 nsew signal output
rlabel metal2 s 75090 119200 75146 120000 6 o[81]
port 367 nsew signal output
rlabel metal2 s 76010 119200 76066 120000 6 o[82]
port 368 nsew signal output
rlabel metal2 s 76930 119200 76986 120000 6 o[83]
port 369 nsew signal output
rlabel metal2 s 77850 119200 77906 120000 6 o[84]
port 370 nsew signal output
rlabel metal2 s 78770 119200 78826 120000 6 o[85]
port 371 nsew signal output
rlabel metal2 s 79690 119200 79746 120000 6 o[86]
port 372 nsew signal output
rlabel metal2 s 80610 119200 80666 120000 6 o[87]
port 373 nsew signal output
rlabel metal2 s 81530 119200 81586 120000 6 o[88]
port 374 nsew signal output
rlabel metal2 s 82450 119200 82506 120000 6 o[89]
port 375 nsew signal output
rlabel metal2 s 7930 119200 7986 120000 6 o[8]
port 376 nsew signal output
rlabel metal2 s 83370 119200 83426 120000 6 o[90]
port 377 nsew signal output
rlabel metal2 s 84290 119200 84346 120000 6 o[91]
port 378 nsew signal output
rlabel metal2 s 85210 119200 85266 120000 6 o[92]
port 379 nsew signal output
rlabel metal2 s 86130 119200 86186 120000 6 o[93]
port 380 nsew signal output
rlabel metal2 s 87050 119200 87106 120000 6 o[94]
port 381 nsew signal output
rlabel metal2 s 87970 119200 88026 120000 6 o[95]
port 382 nsew signal output
rlabel metal2 s 88890 119200 88946 120000 6 o[96]
port 383 nsew signal output
rlabel metal2 s 89810 119200 89866 120000 6 o[97]
port 384 nsew signal output
rlabel metal2 s 90730 119200 90786 120000 6 o[98]
port 385 nsew signal output
rlabel metal2 s 91650 119200 91706 120000 6 o[99]
port 386 nsew signal output
rlabel metal2 s 8850 119200 8906 120000 6 o[9]
port 387 nsew signal output
rlabel metal2 s 118330 119200 118386 120000 6 rst
port 388 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 36087342
string GDS_FILE /scratch/mpw7/caravel_user_project/openlane/multiply_add_64x64/runs/22_07_11_21_36/results/signoff/multiply_add_64x64.magic.gds
string GDS_START 294824
<< end >>

