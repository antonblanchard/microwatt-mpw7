magic
tech sky130A
magscale 1 2
timestamp 1670226251
<< obsli1 >>
rect 1104 2159 108836 107729
<< obsm1 >>
rect 198 1844 110000 107760
<< metal2 >>
rect 1950 109200 2006 110000
rect 2778 109200 2834 110000
rect 3606 109200 3662 110000
rect 4434 109200 4490 110000
rect 5262 109200 5318 110000
rect 6090 109200 6146 110000
rect 6918 109200 6974 110000
rect 7746 109200 7802 110000
rect 8574 109200 8630 110000
rect 9402 109200 9458 110000
rect 10230 109200 10286 110000
rect 11058 109200 11114 110000
rect 11886 109200 11942 110000
rect 12714 109200 12770 110000
rect 13542 109200 13598 110000
rect 14370 109200 14426 110000
rect 15198 109200 15254 110000
rect 16026 109200 16082 110000
rect 16854 109200 16910 110000
rect 17682 109200 17738 110000
rect 18510 109200 18566 110000
rect 19338 109200 19394 110000
rect 20166 109200 20222 110000
rect 20994 109200 21050 110000
rect 21822 109200 21878 110000
rect 22650 109200 22706 110000
rect 23478 109200 23534 110000
rect 24306 109200 24362 110000
rect 25134 109200 25190 110000
rect 25962 109200 26018 110000
rect 26790 109200 26846 110000
rect 27618 109200 27674 110000
rect 28446 109200 28502 110000
rect 29274 109200 29330 110000
rect 30102 109200 30158 110000
rect 30930 109200 30986 110000
rect 31758 109200 31814 110000
rect 32586 109200 32642 110000
rect 33414 109200 33470 110000
rect 34242 109200 34298 110000
rect 35070 109200 35126 110000
rect 35898 109200 35954 110000
rect 36726 109200 36782 110000
rect 37554 109200 37610 110000
rect 38382 109200 38438 110000
rect 39210 109200 39266 110000
rect 40038 109200 40094 110000
rect 40866 109200 40922 110000
rect 41694 109200 41750 110000
rect 42522 109200 42578 110000
rect 43350 109200 43406 110000
rect 44178 109200 44234 110000
rect 45006 109200 45062 110000
rect 45834 109200 45890 110000
rect 46662 109200 46718 110000
rect 47490 109200 47546 110000
rect 48318 109200 48374 110000
rect 49146 109200 49202 110000
rect 49974 109200 50030 110000
rect 50802 109200 50858 110000
rect 51630 109200 51686 110000
rect 52458 109200 52514 110000
rect 53286 109200 53342 110000
rect 54114 109200 54170 110000
rect 54942 109200 54998 110000
rect 55770 109200 55826 110000
rect 56598 109200 56654 110000
rect 57426 109200 57482 110000
rect 58254 109200 58310 110000
rect 59082 109200 59138 110000
rect 59910 109200 59966 110000
rect 60738 109200 60794 110000
rect 61566 109200 61622 110000
rect 62394 109200 62450 110000
rect 63222 109200 63278 110000
rect 64050 109200 64106 110000
rect 64878 109200 64934 110000
rect 65706 109200 65762 110000
rect 66534 109200 66590 110000
rect 67362 109200 67418 110000
rect 68190 109200 68246 110000
rect 69018 109200 69074 110000
rect 69846 109200 69902 110000
rect 70674 109200 70730 110000
rect 71502 109200 71558 110000
rect 72330 109200 72386 110000
rect 73158 109200 73214 110000
rect 73986 109200 74042 110000
rect 74814 109200 74870 110000
rect 75642 109200 75698 110000
rect 76470 109200 76526 110000
rect 77298 109200 77354 110000
rect 78126 109200 78182 110000
rect 78954 109200 79010 110000
rect 79782 109200 79838 110000
rect 80610 109200 80666 110000
rect 81438 109200 81494 110000
rect 82266 109200 82322 110000
rect 83094 109200 83150 110000
rect 83922 109200 83978 110000
rect 84750 109200 84806 110000
rect 85578 109200 85634 110000
rect 86406 109200 86462 110000
rect 87234 109200 87290 110000
rect 88062 109200 88118 110000
rect 88890 109200 88946 110000
rect 89718 109200 89774 110000
rect 90546 109200 90602 110000
rect 91374 109200 91430 110000
rect 92202 109200 92258 110000
rect 93030 109200 93086 110000
rect 93858 109200 93914 110000
rect 94686 109200 94742 110000
rect 95514 109200 95570 110000
rect 96342 109200 96398 110000
rect 97170 109200 97226 110000
rect 97998 109200 98054 110000
rect 98826 109200 98882 110000
rect 99654 109200 99710 110000
rect 100482 109200 100538 110000
rect 101310 109200 101366 110000
rect 102138 109200 102194 110000
rect 102966 109200 103022 110000
rect 103794 109200 103850 110000
rect 104622 109200 104678 110000
rect 105450 109200 105506 110000
rect 106278 109200 106334 110000
rect 107106 109200 107162 110000
rect 107934 109200 107990 110000
rect 2410 0 2466 800
rect 3238 0 3294 800
rect 4066 0 4122 800
rect 4894 0 4950 800
rect 5722 0 5778 800
rect 6550 0 6606 800
rect 7378 0 7434 800
rect 8206 0 8262 800
rect 9034 0 9090 800
rect 9862 0 9918 800
rect 10690 0 10746 800
rect 11518 0 11574 800
rect 12346 0 12402 800
rect 13174 0 13230 800
rect 14002 0 14058 800
rect 14830 0 14886 800
rect 15658 0 15714 800
rect 16486 0 16542 800
rect 17314 0 17370 800
rect 18142 0 18198 800
rect 18970 0 19026 800
rect 19798 0 19854 800
rect 20626 0 20682 800
rect 21454 0 21510 800
rect 22282 0 22338 800
rect 23110 0 23166 800
rect 23938 0 23994 800
rect 24766 0 24822 800
rect 25594 0 25650 800
rect 26422 0 26478 800
rect 27250 0 27306 800
rect 28078 0 28134 800
rect 28906 0 28962 800
rect 29734 0 29790 800
rect 30562 0 30618 800
rect 31390 0 31446 800
rect 32218 0 32274 800
rect 33046 0 33102 800
rect 33874 0 33930 800
rect 34702 0 34758 800
rect 35530 0 35586 800
rect 36358 0 36414 800
rect 37186 0 37242 800
rect 38014 0 38070 800
rect 38842 0 38898 800
rect 39670 0 39726 800
rect 40498 0 40554 800
rect 41326 0 41382 800
rect 42154 0 42210 800
rect 42982 0 43038 800
rect 43810 0 43866 800
rect 44638 0 44694 800
rect 45466 0 45522 800
rect 46294 0 46350 800
rect 47122 0 47178 800
rect 47950 0 48006 800
rect 48778 0 48834 800
rect 49606 0 49662 800
rect 50434 0 50490 800
rect 51262 0 51318 800
rect 52090 0 52146 800
rect 52918 0 52974 800
rect 53746 0 53802 800
rect 54574 0 54630 800
rect 55402 0 55458 800
rect 56230 0 56286 800
rect 57058 0 57114 800
rect 57886 0 57942 800
rect 58714 0 58770 800
rect 59542 0 59598 800
rect 60370 0 60426 800
rect 61198 0 61254 800
rect 62026 0 62082 800
rect 62854 0 62910 800
rect 63682 0 63738 800
rect 64510 0 64566 800
rect 65338 0 65394 800
rect 66166 0 66222 800
rect 66994 0 67050 800
rect 67822 0 67878 800
rect 68650 0 68706 800
rect 69478 0 69534 800
rect 70306 0 70362 800
rect 71134 0 71190 800
rect 71962 0 72018 800
rect 72790 0 72846 800
rect 73618 0 73674 800
rect 74446 0 74502 800
rect 75274 0 75330 800
rect 76102 0 76158 800
rect 76930 0 76986 800
rect 77758 0 77814 800
rect 78586 0 78642 800
rect 79414 0 79470 800
rect 80242 0 80298 800
rect 81070 0 81126 800
rect 81898 0 81954 800
rect 82726 0 82782 800
rect 83554 0 83610 800
rect 84382 0 84438 800
rect 85210 0 85266 800
rect 86038 0 86094 800
rect 86866 0 86922 800
rect 87694 0 87750 800
rect 88522 0 88578 800
rect 89350 0 89406 800
rect 90178 0 90234 800
rect 91006 0 91062 800
rect 91834 0 91890 800
rect 92662 0 92718 800
rect 93490 0 93546 800
rect 94318 0 94374 800
rect 95146 0 95202 800
rect 95974 0 96030 800
rect 96802 0 96858 800
rect 97630 0 97686 800
rect 98458 0 98514 800
rect 99286 0 99342 800
rect 100114 0 100170 800
rect 100942 0 100998 800
rect 101770 0 101826 800
rect 102598 0 102654 800
rect 103426 0 103482 800
rect 104254 0 104310 800
rect 105082 0 105138 800
rect 105910 0 105966 800
rect 106738 0 106794 800
rect 107566 0 107622 800
<< obsm2 >>
rect 124 109144 1894 109290
rect 2062 109144 2722 109290
rect 2890 109144 3550 109290
rect 3718 109144 4378 109290
rect 4546 109144 5206 109290
rect 5374 109144 6034 109290
rect 6202 109144 6862 109290
rect 7030 109144 7690 109290
rect 7858 109144 8518 109290
rect 8686 109144 9346 109290
rect 9514 109144 10174 109290
rect 10342 109144 11002 109290
rect 11170 109144 11830 109290
rect 11998 109144 12658 109290
rect 12826 109144 13486 109290
rect 13654 109144 14314 109290
rect 14482 109144 15142 109290
rect 15310 109144 15970 109290
rect 16138 109144 16798 109290
rect 16966 109144 17626 109290
rect 17794 109144 18454 109290
rect 18622 109144 19282 109290
rect 19450 109144 20110 109290
rect 20278 109144 20938 109290
rect 21106 109144 21766 109290
rect 21934 109144 22594 109290
rect 22762 109144 23422 109290
rect 23590 109144 24250 109290
rect 24418 109144 25078 109290
rect 25246 109144 25906 109290
rect 26074 109144 26734 109290
rect 26902 109144 27562 109290
rect 27730 109144 28390 109290
rect 28558 109144 29218 109290
rect 29386 109144 30046 109290
rect 30214 109144 30874 109290
rect 31042 109144 31702 109290
rect 31870 109144 32530 109290
rect 32698 109144 33358 109290
rect 33526 109144 34186 109290
rect 34354 109144 35014 109290
rect 35182 109144 35842 109290
rect 36010 109144 36670 109290
rect 36838 109144 37498 109290
rect 37666 109144 38326 109290
rect 38494 109144 39154 109290
rect 39322 109144 39982 109290
rect 40150 109144 40810 109290
rect 40978 109144 41638 109290
rect 41806 109144 42466 109290
rect 42634 109144 43294 109290
rect 43462 109144 44122 109290
rect 44290 109144 44950 109290
rect 45118 109144 45778 109290
rect 45946 109144 46606 109290
rect 46774 109144 47434 109290
rect 47602 109144 48262 109290
rect 48430 109144 49090 109290
rect 49258 109144 49918 109290
rect 50086 109144 50746 109290
rect 50914 109144 51574 109290
rect 51742 109144 52402 109290
rect 52570 109144 53230 109290
rect 53398 109144 54058 109290
rect 54226 109144 54886 109290
rect 55054 109144 55714 109290
rect 55882 109144 56542 109290
rect 56710 109144 57370 109290
rect 57538 109144 58198 109290
rect 58366 109144 59026 109290
rect 59194 109144 59854 109290
rect 60022 109144 60682 109290
rect 60850 109144 61510 109290
rect 61678 109144 62338 109290
rect 62506 109144 63166 109290
rect 63334 109144 63994 109290
rect 64162 109144 64822 109290
rect 64990 109144 65650 109290
rect 65818 109144 66478 109290
rect 66646 109144 67306 109290
rect 67474 109144 68134 109290
rect 68302 109144 68962 109290
rect 69130 109144 69790 109290
rect 69958 109144 70618 109290
rect 70786 109144 71446 109290
rect 71614 109144 72274 109290
rect 72442 109144 73102 109290
rect 73270 109144 73930 109290
rect 74098 109144 74758 109290
rect 74926 109144 75586 109290
rect 75754 109144 76414 109290
rect 76582 109144 77242 109290
rect 77410 109144 78070 109290
rect 78238 109144 78898 109290
rect 79066 109144 79726 109290
rect 79894 109144 80554 109290
rect 80722 109144 81382 109290
rect 81550 109144 82210 109290
rect 82378 109144 83038 109290
rect 83206 109144 83866 109290
rect 84034 109144 84694 109290
rect 84862 109144 85522 109290
rect 85690 109144 86350 109290
rect 86518 109144 87178 109290
rect 87346 109144 88006 109290
rect 88174 109144 88834 109290
rect 89002 109144 89662 109290
rect 89830 109144 90490 109290
rect 90658 109144 91318 109290
rect 91486 109144 92146 109290
rect 92314 109144 92974 109290
rect 93142 109144 93802 109290
rect 93970 109144 94630 109290
rect 94798 109144 95458 109290
rect 95626 109144 96286 109290
rect 96454 109144 97114 109290
rect 97282 109144 97942 109290
rect 98110 109144 98770 109290
rect 98938 109144 99598 109290
rect 99766 109144 100426 109290
rect 100594 109144 101254 109290
rect 101422 109144 102082 109290
rect 102250 109144 102910 109290
rect 103078 109144 103738 109290
rect 103906 109144 104566 109290
rect 104734 109144 105394 109290
rect 105562 109144 106222 109290
rect 106390 109144 107050 109290
rect 107218 109144 107878 109290
rect 108046 109144 110000 109290
rect 124 856 110000 109144
rect 124 800 2354 856
rect 2522 800 3182 856
rect 3350 800 4010 856
rect 4178 800 4838 856
rect 5006 800 5666 856
rect 5834 800 6494 856
rect 6662 800 7322 856
rect 7490 800 8150 856
rect 8318 800 8978 856
rect 9146 800 9806 856
rect 9974 800 10634 856
rect 10802 800 11462 856
rect 11630 800 12290 856
rect 12458 800 13118 856
rect 13286 800 13946 856
rect 14114 800 14774 856
rect 14942 800 15602 856
rect 15770 800 16430 856
rect 16598 800 17258 856
rect 17426 800 18086 856
rect 18254 800 18914 856
rect 19082 800 19742 856
rect 19910 800 20570 856
rect 20738 800 21398 856
rect 21566 800 22226 856
rect 22394 800 23054 856
rect 23222 800 23882 856
rect 24050 800 24710 856
rect 24878 800 25538 856
rect 25706 800 26366 856
rect 26534 800 27194 856
rect 27362 800 28022 856
rect 28190 800 28850 856
rect 29018 800 29678 856
rect 29846 800 30506 856
rect 30674 800 31334 856
rect 31502 800 32162 856
rect 32330 800 32990 856
rect 33158 800 33818 856
rect 33986 800 34646 856
rect 34814 800 35474 856
rect 35642 800 36302 856
rect 36470 800 37130 856
rect 37298 800 37958 856
rect 38126 800 38786 856
rect 38954 800 39614 856
rect 39782 800 40442 856
rect 40610 800 41270 856
rect 41438 800 42098 856
rect 42266 800 42926 856
rect 43094 800 43754 856
rect 43922 800 44582 856
rect 44750 800 45410 856
rect 45578 800 46238 856
rect 46406 800 47066 856
rect 47234 800 47894 856
rect 48062 800 48722 856
rect 48890 800 49550 856
rect 49718 800 50378 856
rect 50546 800 51206 856
rect 51374 800 52034 856
rect 52202 800 52862 856
rect 53030 800 53690 856
rect 53858 800 54518 856
rect 54686 800 55346 856
rect 55514 800 56174 856
rect 56342 800 57002 856
rect 57170 800 57830 856
rect 57998 800 58658 856
rect 58826 800 59486 856
rect 59654 800 60314 856
rect 60482 800 61142 856
rect 61310 800 61970 856
rect 62138 800 62798 856
rect 62966 800 63626 856
rect 63794 800 64454 856
rect 64622 800 65282 856
rect 65450 800 66110 856
rect 66278 800 66938 856
rect 67106 800 67766 856
rect 67934 800 68594 856
rect 68762 800 69422 856
rect 69590 800 70250 856
rect 70418 800 71078 856
rect 71246 800 71906 856
rect 72074 800 72734 856
rect 72902 800 73562 856
rect 73730 800 74390 856
rect 74558 800 75218 856
rect 75386 800 76046 856
rect 76214 800 76874 856
rect 77042 800 77702 856
rect 77870 800 78530 856
rect 78698 800 79358 856
rect 79526 800 80186 856
rect 80354 800 81014 856
rect 81182 800 81842 856
rect 82010 800 82670 856
rect 82838 800 83498 856
rect 83666 800 84326 856
rect 84494 800 85154 856
rect 85322 800 85982 856
rect 86150 800 86810 856
rect 86978 800 87638 856
rect 87806 800 88466 856
rect 88634 800 89294 856
rect 89462 800 90122 856
rect 90290 800 90950 856
rect 91118 800 91778 856
rect 91946 800 92606 856
rect 92774 800 93434 856
rect 93602 800 94262 856
rect 94430 800 95090 856
rect 95258 800 95918 856
rect 96086 800 96746 856
rect 96914 800 97574 856
rect 97742 800 98402 856
rect 98570 800 99230 856
rect 99398 800 100058 856
rect 100226 800 100886 856
rect 101054 800 101714 856
rect 101882 800 102542 856
rect 102710 800 103370 856
rect 103538 800 104198 856
rect 104366 800 105026 856
rect 105194 800 105854 856
rect 106022 800 106682 856
rect 106850 800 107510 856
rect 107678 800 110000 856
<< metal3 >>
rect 109200 107176 110000 107296
rect 109200 106360 110000 106480
rect 109200 105544 110000 105664
rect 109200 104728 110000 104848
rect 109200 103912 110000 104032
rect 109200 103096 110000 103216
rect 109200 102280 110000 102400
rect 109200 101464 110000 101584
rect 109200 100648 110000 100768
rect 109200 99832 110000 99952
rect 109200 99016 110000 99136
rect 109200 98200 110000 98320
rect 109200 97384 110000 97504
rect 109200 96568 110000 96688
rect 109200 95752 110000 95872
rect 109200 94936 110000 95056
rect 109200 94120 110000 94240
rect 109200 93304 110000 93424
rect 109200 92488 110000 92608
rect 109200 91672 110000 91792
rect 109200 90856 110000 90976
rect 109200 90040 110000 90160
rect 109200 89224 110000 89344
rect 109200 88408 110000 88528
rect 109200 87592 110000 87712
rect 109200 86776 110000 86896
rect 109200 85960 110000 86080
rect 109200 85144 110000 85264
rect 109200 84328 110000 84448
rect 109200 83512 110000 83632
rect 109200 82696 110000 82816
rect 109200 81880 110000 82000
rect 109200 81064 110000 81184
rect 109200 80248 110000 80368
rect 109200 79432 110000 79552
rect 109200 78616 110000 78736
rect 109200 77800 110000 77920
rect 109200 76984 110000 77104
rect 109200 76168 110000 76288
rect 109200 75352 110000 75472
rect 109200 74536 110000 74656
rect 109200 73720 110000 73840
rect 109200 72904 110000 73024
rect 109200 72088 110000 72208
rect 109200 71272 110000 71392
rect 109200 70456 110000 70576
rect 109200 69640 110000 69760
rect 109200 68824 110000 68944
rect 109200 68008 110000 68128
rect 109200 67192 110000 67312
rect 109200 66376 110000 66496
rect 109200 65560 110000 65680
rect 109200 64744 110000 64864
rect 109200 63928 110000 64048
rect 109200 63112 110000 63232
rect 109200 62296 110000 62416
rect 109200 61480 110000 61600
rect 109200 60664 110000 60784
rect 109200 59848 110000 59968
rect 109200 59032 110000 59152
rect 109200 58216 110000 58336
rect 109200 57400 110000 57520
rect 109200 56584 110000 56704
rect 109200 55768 110000 55888
rect 109200 54952 110000 55072
rect 109200 54136 110000 54256
rect 109200 53320 110000 53440
rect 109200 52504 110000 52624
rect 109200 51688 110000 51808
rect 109200 50872 110000 50992
rect 109200 50056 110000 50176
rect 109200 49240 110000 49360
rect 109200 48424 110000 48544
rect 109200 47608 110000 47728
rect 109200 46792 110000 46912
rect 109200 45976 110000 46096
rect 109200 45160 110000 45280
rect 109200 44344 110000 44464
rect 109200 43528 110000 43648
rect 109200 42712 110000 42832
rect 109200 41896 110000 42016
rect 109200 41080 110000 41200
rect 109200 40264 110000 40384
rect 109200 39448 110000 39568
rect 109200 38632 110000 38752
rect 109200 37816 110000 37936
rect 109200 37000 110000 37120
rect 109200 36184 110000 36304
rect 109200 35368 110000 35488
rect 109200 34552 110000 34672
rect 109200 33736 110000 33856
rect 109200 32920 110000 33040
rect 109200 32104 110000 32224
rect 109200 31288 110000 31408
rect 109200 30472 110000 30592
rect 109200 29656 110000 29776
rect 109200 28840 110000 28960
rect 109200 28024 110000 28144
rect 109200 27208 110000 27328
rect 109200 26392 110000 26512
rect 109200 25576 110000 25696
rect 109200 24760 110000 24880
rect 109200 23944 110000 24064
rect 109200 23128 110000 23248
rect 109200 22312 110000 22432
rect 109200 21496 110000 21616
rect 109200 20680 110000 20800
rect 109200 19864 110000 19984
rect 109200 19048 110000 19168
rect 109200 18232 110000 18352
rect 109200 17416 110000 17536
rect 109200 16600 110000 16720
rect 109200 15784 110000 15904
rect 109200 14968 110000 15088
rect 109200 14152 110000 14272
rect 109200 13336 110000 13456
rect 109200 12520 110000 12640
rect 109200 11704 110000 11824
rect 109200 10888 110000 11008
rect 109200 10072 110000 10192
rect 109200 9256 110000 9376
rect 109200 8440 110000 8560
rect 109200 7624 110000 7744
rect 109200 6808 110000 6928
rect 109200 5992 110000 6112
rect 109200 5176 110000 5296
rect 109200 4360 110000 4480
rect 109200 3544 110000 3664
rect 109200 2728 110000 2848
<< obsm3 >>
rect 381 107376 109927 107745
rect 381 107096 109120 107376
rect 381 106560 109927 107096
rect 381 106280 109120 106560
rect 381 105744 109927 106280
rect 381 105464 109120 105744
rect 381 104928 109927 105464
rect 381 104648 109120 104928
rect 381 104112 109927 104648
rect 381 103832 109120 104112
rect 381 103296 109927 103832
rect 381 103016 109120 103296
rect 381 102480 109927 103016
rect 381 102200 109120 102480
rect 381 101664 109927 102200
rect 381 101384 109120 101664
rect 381 100848 109927 101384
rect 381 100568 109120 100848
rect 381 100032 109927 100568
rect 381 99752 109120 100032
rect 381 99216 109927 99752
rect 381 98936 109120 99216
rect 381 98400 109927 98936
rect 381 98120 109120 98400
rect 381 97584 109927 98120
rect 381 97304 109120 97584
rect 381 96768 109927 97304
rect 381 96488 109120 96768
rect 381 95952 109927 96488
rect 381 95672 109120 95952
rect 381 95136 109927 95672
rect 381 94856 109120 95136
rect 381 94320 109927 94856
rect 381 94040 109120 94320
rect 381 93504 109927 94040
rect 381 93224 109120 93504
rect 381 92688 109927 93224
rect 381 92408 109120 92688
rect 381 91872 109927 92408
rect 381 91592 109120 91872
rect 381 91056 109927 91592
rect 381 90776 109120 91056
rect 381 90240 109927 90776
rect 381 89960 109120 90240
rect 381 89424 109927 89960
rect 381 89144 109120 89424
rect 381 88608 109927 89144
rect 381 88328 109120 88608
rect 381 87792 109927 88328
rect 381 87512 109120 87792
rect 381 86976 109927 87512
rect 381 86696 109120 86976
rect 381 86160 109927 86696
rect 381 85880 109120 86160
rect 381 85344 109927 85880
rect 381 85064 109120 85344
rect 381 84528 109927 85064
rect 381 84248 109120 84528
rect 381 83712 109927 84248
rect 381 83432 109120 83712
rect 381 82896 109927 83432
rect 381 82616 109120 82896
rect 381 82080 109927 82616
rect 381 81800 109120 82080
rect 381 81264 109927 81800
rect 381 80984 109120 81264
rect 381 80448 109927 80984
rect 381 80168 109120 80448
rect 381 79632 109927 80168
rect 381 79352 109120 79632
rect 381 78816 109927 79352
rect 381 78536 109120 78816
rect 381 78000 109927 78536
rect 381 77720 109120 78000
rect 381 77184 109927 77720
rect 381 76904 109120 77184
rect 381 76368 109927 76904
rect 381 76088 109120 76368
rect 381 75552 109927 76088
rect 381 75272 109120 75552
rect 381 74736 109927 75272
rect 381 74456 109120 74736
rect 381 73920 109927 74456
rect 381 73640 109120 73920
rect 381 73104 109927 73640
rect 381 72824 109120 73104
rect 381 72288 109927 72824
rect 381 72008 109120 72288
rect 381 71472 109927 72008
rect 381 71192 109120 71472
rect 381 70656 109927 71192
rect 381 70376 109120 70656
rect 381 69840 109927 70376
rect 381 69560 109120 69840
rect 381 69024 109927 69560
rect 381 68744 109120 69024
rect 381 68208 109927 68744
rect 381 67928 109120 68208
rect 381 67392 109927 67928
rect 381 67112 109120 67392
rect 381 66576 109927 67112
rect 381 66296 109120 66576
rect 381 65760 109927 66296
rect 381 65480 109120 65760
rect 381 64944 109927 65480
rect 381 64664 109120 64944
rect 381 64128 109927 64664
rect 381 63848 109120 64128
rect 381 63312 109927 63848
rect 381 63032 109120 63312
rect 381 62496 109927 63032
rect 381 62216 109120 62496
rect 381 61680 109927 62216
rect 381 61400 109120 61680
rect 381 60864 109927 61400
rect 381 60584 109120 60864
rect 381 60048 109927 60584
rect 381 59768 109120 60048
rect 381 59232 109927 59768
rect 381 58952 109120 59232
rect 381 58416 109927 58952
rect 381 58136 109120 58416
rect 381 57600 109927 58136
rect 381 57320 109120 57600
rect 381 56784 109927 57320
rect 381 56504 109120 56784
rect 381 55968 109927 56504
rect 381 55688 109120 55968
rect 381 55152 109927 55688
rect 381 54872 109120 55152
rect 381 54336 109927 54872
rect 381 54056 109120 54336
rect 381 53520 109927 54056
rect 381 53240 109120 53520
rect 381 52704 109927 53240
rect 381 52424 109120 52704
rect 381 51888 109927 52424
rect 381 51608 109120 51888
rect 381 51072 109927 51608
rect 381 50792 109120 51072
rect 381 50256 109927 50792
rect 381 49976 109120 50256
rect 381 49440 109927 49976
rect 381 49160 109120 49440
rect 381 48624 109927 49160
rect 381 48344 109120 48624
rect 381 47808 109927 48344
rect 381 47528 109120 47808
rect 381 46992 109927 47528
rect 381 46712 109120 46992
rect 381 46176 109927 46712
rect 381 45896 109120 46176
rect 381 45360 109927 45896
rect 381 45080 109120 45360
rect 381 44544 109927 45080
rect 381 44264 109120 44544
rect 381 43728 109927 44264
rect 381 43448 109120 43728
rect 381 42912 109927 43448
rect 381 42632 109120 42912
rect 381 42096 109927 42632
rect 381 41816 109120 42096
rect 381 41280 109927 41816
rect 381 41000 109120 41280
rect 381 40464 109927 41000
rect 381 40184 109120 40464
rect 381 39648 109927 40184
rect 381 39368 109120 39648
rect 381 38832 109927 39368
rect 381 38552 109120 38832
rect 381 38016 109927 38552
rect 381 37736 109120 38016
rect 381 37200 109927 37736
rect 381 36920 109120 37200
rect 381 36384 109927 36920
rect 381 36104 109120 36384
rect 381 35568 109927 36104
rect 381 35288 109120 35568
rect 381 34752 109927 35288
rect 381 34472 109120 34752
rect 381 33936 109927 34472
rect 381 33656 109120 33936
rect 381 33120 109927 33656
rect 381 32840 109120 33120
rect 381 32304 109927 32840
rect 381 32024 109120 32304
rect 381 31488 109927 32024
rect 381 31208 109120 31488
rect 381 30672 109927 31208
rect 381 30392 109120 30672
rect 381 29856 109927 30392
rect 381 29576 109120 29856
rect 381 29040 109927 29576
rect 381 28760 109120 29040
rect 381 28224 109927 28760
rect 381 27944 109120 28224
rect 381 27408 109927 27944
rect 381 27128 109120 27408
rect 381 26592 109927 27128
rect 381 26312 109120 26592
rect 381 25776 109927 26312
rect 381 25496 109120 25776
rect 381 24960 109927 25496
rect 381 24680 109120 24960
rect 381 24144 109927 24680
rect 381 23864 109120 24144
rect 381 23328 109927 23864
rect 381 23048 109120 23328
rect 381 22512 109927 23048
rect 381 22232 109120 22512
rect 381 21696 109927 22232
rect 381 21416 109120 21696
rect 381 20880 109927 21416
rect 381 20600 109120 20880
rect 381 20064 109927 20600
rect 381 19784 109120 20064
rect 381 19248 109927 19784
rect 381 18968 109120 19248
rect 381 18432 109927 18968
rect 381 18152 109120 18432
rect 381 17616 109927 18152
rect 381 17336 109120 17616
rect 381 16800 109927 17336
rect 381 16520 109120 16800
rect 381 15984 109927 16520
rect 381 15704 109120 15984
rect 381 15168 109927 15704
rect 381 14888 109120 15168
rect 381 14352 109927 14888
rect 381 14072 109120 14352
rect 381 13536 109927 14072
rect 381 13256 109120 13536
rect 381 12720 109927 13256
rect 381 12440 109120 12720
rect 381 11904 109927 12440
rect 381 11624 109120 11904
rect 381 11088 109927 11624
rect 381 10808 109120 11088
rect 381 10272 109927 10808
rect 381 9992 109120 10272
rect 381 9456 109927 9992
rect 381 9176 109120 9456
rect 381 8640 109927 9176
rect 381 8360 109120 8640
rect 381 7824 109927 8360
rect 381 7544 109120 7824
rect 381 7008 109927 7544
rect 381 6728 109120 7008
rect 381 6192 109927 6728
rect 381 5912 109120 6192
rect 381 5376 109927 5912
rect 381 5096 109120 5376
rect 381 4560 109927 5096
rect 381 4280 109120 4560
rect 381 3744 109927 4280
rect 381 3464 109120 3744
rect 381 2928 109927 3464
rect 381 2648 109120 2928
rect 381 2143 109927 2648
<< metal4 >>
rect 1794 2128 2414 107760
rect 19794 2128 20414 107760
rect 37794 2128 38414 107760
rect 55794 2128 56414 107760
rect 73794 2128 74414 107760
rect 91794 2128 92414 107760
<< obsm4 >>
rect 427 2619 1714 107269
rect 2494 2619 19714 107269
rect 20494 2619 37714 107269
rect 38494 2619 55714 107269
rect 56494 2619 73714 107269
rect 74494 2619 91714 107269
rect 92494 2619 109421 107269
<< labels >>
rlabel metal4 s 19794 2128 20414 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 55794 2128 56414 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 91794 2128 92414 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1794 2128 2414 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 37794 2128 38414 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 73794 2128 74414 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 109200 3544 110000 3664 6 a[0]
port 3 nsew signal input
rlabel metal3 s 109200 11704 110000 11824 6 a[10]
port 4 nsew signal input
rlabel metal3 s 109200 12520 110000 12640 6 a[11]
port 5 nsew signal input
rlabel metal3 s 109200 13336 110000 13456 6 a[12]
port 6 nsew signal input
rlabel metal3 s 109200 14152 110000 14272 6 a[13]
port 7 nsew signal input
rlabel metal3 s 109200 14968 110000 15088 6 a[14]
port 8 nsew signal input
rlabel metal3 s 109200 15784 110000 15904 6 a[15]
port 9 nsew signal input
rlabel metal3 s 109200 16600 110000 16720 6 a[16]
port 10 nsew signal input
rlabel metal3 s 109200 17416 110000 17536 6 a[17]
port 11 nsew signal input
rlabel metal3 s 109200 18232 110000 18352 6 a[18]
port 12 nsew signal input
rlabel metal3 s 109200 19048 110000 19168 6 a[19]
port 13 nsew signal input
rlabel metal3 s 109200 4360 110000 4480 6 a[1]
port 14 nsew signal input
rlabel metal3 s 109200 19864 110000 19984 6 a[20]
port 15 nsew signal input
rlabel metal3 s 109200 20680 110000 20800 6 a[21]
port 16 nsew signal input
rlabel metal3 s 109200 21496 110000 21616 6 a[22]
port 17 nsew signal input
rlabel metal3 s 109200 22312 110000 22432 6 a[23]
port 18 nsew signal input
rlabel metal3 s 109200 23128 110000 23248 6 a[24]
port 19 nsew signal input
rlabel metal3 s 109200 23944 110000 24064 6 a[25]
port 20 nsew signal input
rlabel metal3 s 109200 24760 110000 24880 6 a[26]
port 21 nsew signal input
rlabel metal3 s 109200 25576 110000 25696 6 a[27]
port 22 nsew signal input
rlabel metal3 s 109200 26392 110000 26512 6 a[28]
port 23 nsew signal input
rlabel metal3 s 109200 27208 110000 27328 6 a[29]
port 24 nsew signal input
rlabel metal3 s 109200 5176 110000 5296 6 a[2]
port 25 nsew signal input
rlabel metal3 s 109200 28024 110000 28144 6 a[30]
port 26 nsew signal input
rlabel metal3 s 109200 28840 110000 28960 6 a[31]
port 27 nsew signal input
rlabel metal3 s 109200 29656 110000 29776 6 a[32]
port 28 nsew signal input
rlabel metal3 s 109200 30472 110000 30592 6 a[33]
port 29 nsew signal input
rlabel metal3 s 109200 31288 110000 31408 6 a[34]
port 30 nsew signal input
rlabel metal3 s 109200 32104 110000 32224 6 a[35]
port 31 nsew signal input
rlabel metal3 s 109200 32920 110000 33040 6 a[36]
port 32 nsew signal input
rlabel metal3 s 109200 33736 110000 33856 6 a[37]
port 33 nsew signal input
rlabel metal3 s 109200 34552 110000 34672 6 a[38]
port 34 nsew signal input
rlabel metal3 s 109200 35368 110000 35488 6 a[39]
port 35 nsew signal input
rlabel metal3 s 109200 5992 110000 6112 6 a[3]
port 36 nsew signal input
rlabel metal3 s 109200 36184 110000 36304 6 a[40]
port 37 nsew signal input
rlabel metal3 s 109200 37000 110000 37120 6 a[41]
port 38 nsew signal input
rlabel metal3 s 109200 37816 110000 37936 6 a[42]
port 39 nsew signal input
rlabel metal3 s 109200 38632 110000 38752 6 a[43]
port 40 nsew signal input
rlabel metal3 s 109200 39448 110000 39568 6 a[44]
port 41 nsew signal input
rlabel metal3 s 109200 40264 110000 40384 6 a[45]
port 42 nsew signal input
rlabel metal3 s 109200 41080 110000 41200 6 a[46]
port 43 nsew signal input
rlabel metal3 s 109200 41896 110000 42016 6 a[47]
port 44 nsew signal input
rlabel metal3 s 109200 42712 110000 42832 6 a[48]
port 45 nsew signal input
rlabel metal3 s 109200 43528 110000 43648 6 a[49]
port 46 nsew signal input
rlabel metal3 s 109200 6808 110000 6928 6 a[4]
port 47 nsew signal input
rlabel metal3 s 109200 44344 110000 44464 6 a[50]
port 48 nsew signal input
rlabel metal3 s 109200 45160 110000 45280 6 a[51]
port 49 nsew signal input
rlabel metal3 s 109200 45976 110000 46096 6 a[52]
port 50 nsew signal input
rlabel metal3 s 109200 46792 110000 46912 6 a[53]
port 51 nsew signal input
rlabel metal3 s 109200 47608 110000 47728 6 a[54]
port 52 nsew signal input
rlabel metal3 s 109200 48424 110000 48544 6 a[55]
port 53 nsew signal input
rlabel metal3 s 109200 49240 110000 49360 6 a[56]
port 54 nsew signal input
rlabel metal3 s 109200 50056 110000 50176 6 a[57]
port 55 nsew signal input
rlabel metal3 s 109200 50872 110000 50992 6 a[58]
port 56 nsew signal input
rlabel metal3 s 109200 51688 110000 51808 6 a[59]
port 57 nsew signal input
rlabel metal3 s 109200 7624 110000 7744 6 a[5]
port 58 nsew signal input
rlabel metal3 s 109200 52504 110000 52624 6 a[60]
port 59 nsew signal input
rlabel metal3 s 109200 53320 110000 53440 6 a[61]
port 60 nsew signal input
rlabel metal3 s 109200 54136 110000 54256 6 a[62]
port 61 nsew signal input
rlabel metal3 s 109200 54952 110000 55072 6 a[63]
port 62 nsew signal input
rlabel metal3 s 109200 8440 110000 8560 6 a[6]
port 63 nsew signal input
rlabel metal3 s 109200 9256 110000 9376 6 a[7]
port 64 nsew signal input
rlabel metal3 s 109200 10072 110000 10192 6 a[8]
port 65 nsew signal input
rlabel metal3 s 109200 10888 110000 11008 6 a[9]
port 66 nsew signal input
rlabel metal3 s 109200 55768 110000 55888 6 b[0]
port 67 nsew signal input
rlabel metal3 s 109200 63928 110000 64048 6 b[10]
port 68 nsew signal input
rlabel metal3 s 109200 64744 110000 64864 6 b[11]
port 69 nsew signal input
rlabel metal3 s 109200 65560 110000 65680 6 b[12]
port 70 nsew signal input
rlabel metal3 s 109200 66376 110000 66496 6 b[13]
port 71 nsew signal input
rlabel metal3 s 109200 67192 110000 67312 6 b[14]
port 72 nsew signal input
rlabel metal3 s 109200 68008 110000 68128 6 b[15]
port 73 nsew signal input
rlabel metal3 s 109200 68824 110000 68944 6 b[16]
port 74 nsew signal input
rlabel metal3 s 109200 69640 110000 69760 6 b[17]
port 75 nsew signal input
rlabel metal3 s 109200 70456 110000 70576 6 b[18]
port 76 nsew signal input
rlabel metal3 s 109200 71272 110000 71392 6 b[19]
port 77 nsew signal input
rlabel metal3 s 109200 56584 110000 56704 6 b[1]
port 78 nsew signal input
rlabel metal3 s 109200 72088 110000 72208 6 b[20]
port 79 nsew signal input
rlabel metal3 s 109200 72904 110000 73024 6 b[21]
port 80 nsew signal input
rlabel metal3 s 109200 73720 110000 73840 6 b[22]
port 81 nsew signal input
rlabel metal3 s 109200 74536 110000 74656 6 b[23]
port 82 nsew signal input
rlabel metal3 s 109200 75352 110000 75472 6 b[24]
port 83 nsew signal input
rlabel metal3 s 109200 76168 110000 76288 6 b[25]
port 84 nsew signal input
rlabel metal3 s 109200 76984 110000 77104 6 b[26]
port 85 nsew signal input
rlabel metal3 s 109200 77800 110000 77920 6 b[27]
port 86 nsew signal input
rlabel metal3 s 109200 78616 110000 78736 6 b[28]
port 87 nsew signal input
rlabel metal3 s 109200 79432 110000 79552 6 b[29]
port 88 nsew signal input
rlabel metal3 s 109200 57400 110000 57520 6 b[2]
port 89 nsew signal input
rlabel metal3 s 109200 80248 110000 80368 6 b[30]
port 90 nsew signal input
rlabel metal3 s 109200 81064 110000 81184 6 b[31]
port 91 nsew signal input
rlabel metal3 s 109200 81880 110000 82000 6 b[32]
port 92 nsew signal input
rlabel metal3 s 109200 82696 110000 82816 6 b[33]
port 93 nsew signal input
rlabel metal3 s 109200 83512 110000 83632 6 b[34]
port 94 nsew signal input
rlabel metal3 s 109200 84328 110000 84448 6 b[35]
port 95 nsew signal input
rlabel metal3 s 109200 85144 110000 85264 6 b[36]
port 96 nsew signal input
rlabel metal3 s 109200 85960 110000 86080 6 b[37]
port 97 nsew signal input
rlabel metal3 s 109200 86776 110000 86896 6 b[38]
port 98 nsew signal input
rlabel metal3 s 109200 87592 110000 87712 6 b[39]
port 99 nsew signal input
rlabel metal3 s 109200 58216 110000 58336 6 b[3]
port 100 nsew signal input
rlabel metal3 s 109200 88408 110000 88528 6 b[40]
port 101 nsew signal input
rlabel metal3 s 109200 89224 110000 89344 6 b[41]
port 102 nsew signal input
rlabel metal3 s 109200 90040 110000 90160 6 b[42]
port 103 nsew signal input
rlabel metal3 s 109200 90856 110000 90976 6 b[43]
port 104 nsew signal input
rlabel metal3 s 109200 91672 110000 91792 6 b[44]
port 105 nsew signal input
rlabel metal3 s 109200 92488 110000 92608 6 b[45]
port 106 nsew signal input
rlabel metal3 s 109200 93304 110000 93424 6 b[46]
port 107 nsew signal input
rlabel metal3 s 109200 94120 110000 94240 6 b[47]
port 108 nsew signal input
rlabel metal3 s 109200 94936 110000 95056 6 b[48]
port 109 nsew signal input
rlabel metal3 s 109200 95752 110000 95872 6 b[49]
port 110 nsew signal input
rlabel metal3 s 109200 59032 110000 59152 6 b[4]
port 111 nsew signal input
rlabel metal3 s 109200 96568 110000 96688 6 b[50]
port 112 nsew signal input
rlabel metal3 s 109200 97384 110000 97504 6 b[51]
port 113 nsew signal input
rlabel metal3 s 109200 98200 110000 98320 6 b[52]
port 114 nsew signal input
rlabel metal3 s 109200 99016 110000 99136 6 b[53]
port 115 nsew signal input
rlabel metal3 s 109200 99832 110000 99952 6 b[54]
port 116 nsew signal input
rlabel metal3 s 109200 100648 110000 100768 6 b[55]
port 117 nsew signal input
rlabel metal3 s 109200 101464 110000 101584 6 b[56]
port 118 nsew signal input
rlabel metal3 s 109200 102280 110000 102400 6 b[57]
port 119 nsew signal input
rlabel metal3 s 109200 103096 110000 103216 6 b[58]
port 120 nsew signal input
rlabel metal3 s 109200 103912 110000 104032 6 b[59]
port 121 nsew signal input
rlabel metal3 s 109200 59848 110000 59968 6 b[5]
port 122 nsew signal input
rlabel metal3 s 109200 104728 110000 104848 6 b[60]
port 123 nsew signal input
rlabel metal3 s 109200 105544 110000 105664 6 b[61]
port 124 nsew signal input
rlabel metal3 s 109200 106360 110000 106480 6 b[62]
port 125 nsew signal input
rlabel metal3 s 109200 107176 110000 107296 6 b[63]
port 126 nsew signal input
rlabel metal3 s 109200 60664 110000 60784 6 b[6]
port 127 nsew signal input
rlabel metal3 s 109200 61480 110000 61600 6 b[7]
port 128 nsew signal input
rlabel metal3 s 109200 62296 110000 62416 6 b[8]
port 129 nsew signal input
rlabel metal3 s 109200 63112 110000 63232 6 b[9]
port 130 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 c[0]
port 131 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 c[100]
port 132 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 c[101]
port 133 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 c[102]
port 134 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 c[103]
port 135 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 c[104]
port 136 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 c[105]
port 137 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 c[106]
port 138 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 c[107]
port 139 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 c[108]
port 140 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 c[109]
port 141 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 c[10]
port 142 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 c[110]
port 143 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 c[111]
port 144 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 c[112]
port 145 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 c[113]
port 146 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 c[114]
port 147 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 c[115]
port 148 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 c[116]
port 149 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 c[117]
port 150 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 c[118]
port 151 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 c[119]
port 152 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 c[11]
port 153 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 c[120]
port 154 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 c[121]
port 155 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 c[122]
port 156 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 c[123]
port 157 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 c[124]
port 158 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 c[125]
port 159 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 c[126]
port 160 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 c[127]
port 161 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 c[12]
port 162 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 c[13]
port 163 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 c[14]
port 164 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 c[15]
port 165 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 c[16]
port 166 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 c[17]
port 167 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 c[18]
port 168 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 c[19]
port 169 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 c[1]
port 170 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 c[20]
port 171 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 c[21]
port 172 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 c[22]
port 173 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 c[23]
port 174 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 c[24]
port 175 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 c[25]
port 176 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 c[26]
port 177 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 c[27]
port 178 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 c[28]
port 179 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 c[29]
port 180 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 c[2]
port 181 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 c[30]
port 182 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 c[31]
port 183 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 c[32]
port 184 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 c[33]
port 185 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 c[34]
port 186 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 c[35]
port 187 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 c[36]
port 188 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 c[37]
port 189 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 c[38]
port 190 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 c[39]
port 191 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 c[3]
port 192 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 c[40]
port 193 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 c[41]
port 194 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 c[42]
port 195 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 c[43]
port 196 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 c[44]
port 197 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 c[45]
port 198 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 c[46]
port 199 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 c[47]
port 200 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 c[48]
port 201 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 c[49]
port 202 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 c[4]
port 203 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 c[50]
port 204 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 c[51]
port 205 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 c[52]
port 206 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 c[53]
port 207 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 c[54]
port 208 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 c[55]
port 209 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 c[56]
port 210 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 c[57]
port 211 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 c[58]
port 212 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 c[59]
port 213 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 c[5]
port 214 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 c[60]
port 215 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 c[61]
port 216 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 c[62]
port 217 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 c[63]
port 218 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 c[64]
port 219 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 c[65]
port 220 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 c[66]
port 221 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 c[67]
port 222 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 c[68]
port 223 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 c[69]
port 224 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 c[6]
port 225 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 c[70]
port 226 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 c[71]
port 227 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 c[72]
port 228 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 c[73]
port 229 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 c[74]
port 230 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 c[75]
port 231 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 c[76]
port 232 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 c[77]
port 233 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 c[78]
port 234 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 c[79]
port 235 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 c[7]
port 236 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 c[80]
port 237 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 c[81]
port 238 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 c[82]
port 239 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 c[83]
port 240 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 c[84]
port 241 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 c[85]
port 242 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 c[86]
port 243 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 c[87]
port 244 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 c[88]
port 245 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 c[89]
port 246 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 c[8]
port 247 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 c[90]
port 248 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 c[91]
port 249 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 c[92]
port 250 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 c[93]
port 251 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 c[94]
port 252 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 c[95]
port 253 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 c[96]
port 254 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 c[97]
port 255 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 c[98]
port 256 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 c[99]
port 257 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 c[9]
port 258 nsew signal input
rlabel metal3 s 109200 2728 110000 2848 6 clk
port 259 nsew signal input
rlabel metal2 s 1950 109200 2006 110000 6 o[0]
port 260 nsew signal output
rlabel metal2 s 84750 109200 84806 110000 6 o[100]
port 261 nsew signal output
rlabel metal2 s 85578 109200 85634 110000 6 o[101]
port 262 nsew signal output
rlabel metal2 s 86406 109200 86462 110000 6 o[102]
port 263 nsew signal output
rlabel metal2 s 87234 109200 87290 110000 6 o[103]
port 264 nsew signal output
rlabel metal2 s 88062 109200 88118 110000 6 o[104]
port 265 nsew signal output
rlabel metal2 s 88890 109200 88946 110000 6 o[105]
port 266 nsew signal output
rlabel metal2 s 89718 109200 89774 110000 6 o[106]
port 267 nsew signal output
rlabel metal2 s 90546 109200 90602 110000 6 o[107]
port 268 nsew signal output
rlabel metal2 s 91374 109200 91430 110000 6 o[108]
port 269 nsew signal output
rlabel metal2 s 92202 109200 92258 110000 6 o[109]
port 270 nsew signal output
rlabel metal2 s 10230 109200 10286 110000 6 o[10]
port 271 nsew signal output
rlabel metal2 s 93030 109200 93086 110000 6 o[110]
port 272 nsew signal output
rlabel metal2 s 93858 109200 93914 110000 6 o[111]
port 273 nsew signal output
rlabel metal2 s 94686 109200 94742 110000 6 o[112]
port 274 nsew signal output
rlabel metal2 s 95514 109200 95570 110000 6 o[113]
port 275 nsew signal output
rlabel metal2 s 96342 109200 96398 110000 6 o[114]
port 276 nsew signal output
rlabel metal2 s 97170 109200 97226 110000 6 o[115]
port 277 nsew signal output
rlabel metal2 s 97998 109200 98054 110000 6 o[116]
port 278 nsew signal output
rlabel metal2 s 98826 109200 98882 110000 6 o[117]
port 279 nsew signal output
rlabel metal2 s 99654 109200 99710 110000 6 o[118]
port 280 nsew signal output
rlabel metal2 s 100482 109200 100538 110000 6 o[119]
port 281 nsew signal output
rlabel metal2 s 11058 109200 11114 110000 6 o[11]
port 282 nsew signal output
rlabel metal2 s 101310 109200 101366 110000 6 o[120]
port 283 nsew signal output
rlabel metal2 s 102138 109200 102194 110000 6 o[121]
port 284 nsew signal output
rlabel metal2 s 102966 109200 103022 110000 6 o[122]
port 285 nsew signal output
rlabel metal2 s 103794 109200 103850 110000 6 o[123]
port 286 nsew signal output
rlabel metal2 s 104622 109200 104678 110000 6 o[124]
port 287 nsew signal output
rlabel metal2 s 105450 109200 105506 110000 6 o[125]
port 288 nsew signal output
rlabel metal2 s 106278 109200 106334 110000 6 o[126]
port 289 nsew signal output
rlabel metal2 s 107106 109200 107162 110000 6 o[127]
port 290 nsew signal output
rlabel metal2 s 11886 109200 11942 110000 6 o[12]
port 291 nsew signal output
rlabel metal2 s 12714 109200 12770 110000 6 o[13]
port 292 nsew signal output
rlabel metal2 s 13542 109200 13598 110000 6 o[14]
port 293 nsew signal output
rlabel metal2 s 14370 109200 14426 110000 6 o[15]
port 294 nsew signal output
rlabel metal2 s 15198 109200 15254 110000 6 o[16]
port 295 nsew signal output
rlabel metal2 s 16026 109200 16082 110000 6 o[17]
port 296 nsew signal output
rlabel metal2 s 16854 109200 16910 110000 6 o[18]
port 297 nsew signal output
rlabel metal2 s 17682 109200 17738 110000 6 o[19]
port 298 nsew signal output
rlabel metal2 s 2778 109200 2834 110000 6 o[1]
port 299 nsew signal output
rlabel metal2 s 18510 109200 18566 110000 6 o[20]
port 300 nsew signal output
rlabel metal2 s 19338 109200 19394 110000 6 o[21]
port 301 nsew signal output
rlabel metal2 s 20166 109200 20222 110000 6 o[22]
port 302 nsew signal output
rlabel metal2 s 20994 109200 21050 110000 6 o[23]
port 303 nsew signal output
rlabel metal2 s 21822 109200 21878 110000 6 o[24]
port 304 nsew signal output
rlabel metal2 s 22650 109200 22706 110000 6 o[25]
port 305 nsew signal output
rlabel metal2 s 23478 109200 23534 110000 6 o[26]
port 306 nsew signal output
rlabel metal2 s 24306 109200 24362 110000 6 o[27]
port 307 nsew signal output
rlabel metal2 s 25134 109200 25190 110000 6 o[28]
port 308 nsew signal output
rlabel metal2 s 25962 109200 26018 110000 6 o[29]
port 309 nsew signal output
rlabel metal2 s 3606 109200 3662 110000 6 o[2]
port 310 nsew signal output
rlabel metal2 s 26790 109200 26846 110000 6 o[30]
port 311 nsew signal output
rlabel metal2 s 27618 109200 27674 110000 6 o[31]
port 312 nsew signal output
rlabel metal2 s 28446 109200 28502 110000 6 o[32]
port 313 nsew signal output
rlabel metal2 s 29274 109200 29330 110000 6 o[33]
port 314 nsew signal output
rlabel metal2 s 30102 109200 30158 110000 6 o[34]
port 315 nsew signal output
rlabel metal2 s 30930 109200 30986 110000 6 o[35]
port 316 nsew signal output
rlabel metal2 s 31758 109200 31814 110000 6 o[36]
port 317 nsew signal output
rlabel metal2 s 32586 109200 32642 110000 6 o[37]
port 318 nsew signal output
rlabel metal2 s 33414 109200 33470 110000 6 o[38]
port 319 nsew signal output
rlabel metal2 s 34242 109200 34298 110000 6 o[39]
port 320 nsew signal output
rlabel metal2 s 4434 109200 4490 110000 6 o[3]
port 321 nsew signal output
rlabel metal2 s 35070 109200 35126 110000 6 o[40]
port 322 nsew signal output
rlabel metal2 s 35898 109200 35954 110000 6 o[41]
port 323 nsew signal output
rlabel metal2 s 36726 109200 36782 110000 6 o[42]
port 324 nsew signal output
rlabel metal2 s 37554 109200 37610 110000 6 o[43]
port 325 nsew signal output
rlabel metal2 s 38382 109200 38438 110000 6 o[44]
port 326 nsew signal output
rlabel metal2 s 39210 109200 39266 110000 6 o[45]
port 327 nsew signal output
rlabel metal2 s 40038 109200 40094 110000 6 o[46]
port 328 nsew signal output
rlabel metal2 s 40866 109200 40922 110000 6 o[47]
port 329 nsew signal output
rlabel metal2 s 41694 109200 41750 110000 6 o[48]
port 330 nsew signal output
rlabel metal2 s 42522 109200 42578 110000 6 o[49]
port 331 nsew signal output
rlabel metal2 s 5262 109200 5318 110000 6 o[4]
port 332 nsew signal output
rlabel metal2 s 43350 109200 43406 110000 6 o[50]
port 333 nsew signal output
rlabel metal2 s 44178 109200 44234 110000 6 o[51]
port 334 nsew signal output
rlabel metal2 s 45006 109200 45062 110000 6 o[52]
port 335 nsew signal output
rlabel metal2 s 45834 109200 45890 110000 6 o[53]
port 336 nsew signal output
rlabel metal2 s 46662 109200 46718 110000 6 o[54]
port 337 nsew signal output
rlabel metal2 s 47490 109200 47546 110000 6 o[55]
port 338 nsew signal output
rlabel metal2 s 48318 109200 48374 110000 6 o[56]
port 339 nsew signal output
rlabel metal2 s 49146 109200 49202 110000 6 o[57]
port 340 nsew signal output
rlabel metal2 s 49974 109200 50030 110000 6 o[58]
port 341 nsew signal output
rlabel metal2 s 50802 109200 50858 110000 6 o[59]
port 342 nsew signal output
rlabel metal2 s 6090 109200 6146 110000 6 o[5]
port 343 nsew signal output
rlabel metal2 s 51630 109200 51686 110000 6 o[60]
port 344 nsew signal output
rlabel metal2 s 52458 109200 52514 110000 6 o[61]
port 345 nsew signal output
rlabel metal2 s 53286 109200 53342 110000 6 o[62]
port 346 nsew signal output
rlabel metal2 s 54114 109200 54170 110000 6 o[63]
port 347 nsew signal output
rlabel metal2 s 54942 109200 54998 110000 6 o[64]
port 348 nsew signal output
rlabel metal2 s 55770 109200 55826 110000 6 o[65]
port 349 nsew signal output
rlabel metal2 s 56598 109200 56654 110000 6 o[66]
port 350 nsew signal output
rlabel metal2 s 57426 109200 57482 110000 6 o[67]
port 351 nsew signal output
rlabel metal2 s 58254 109200 58310 110000 6 o[68]
port 352 nsew signal output
rlabel metal2 s 59082 109200 59138 110000 6 o[69]
port 353 nsew signal output
rlabel metal2 s 6918 109200 6974 110000 6 o[6]
port 354 nsew signal output
rlabel metal2 s 59910 109200 59966 110000 6 o[70]
port 355 nsew signal output
rlabel metal2 s 60738 109200 60794 110000 6 o[71]
port 356 nsew signal output
rlabel metal2 s 61566 109200 61622 110000 6 o[72]
port 357 nsew signal output
rlabel metal2 s 62394 109200 62450 110000 6 o[73]
port 358 nsew signal output
rlabel metal2 s 63222 109200 63278 110000 6 o[74]
port 359 nsew signal output
rlabel metal2 s 64050 109200 64106 110000 6 o[75]
port 360 nsew signal output
rlabel metal2 s 64878 109200 64934 110000 6 o[76]
port 361 nsew signal output
rlabel metal2 s 65706 109200 65762 110000 6 o[77]
port 362 nsew signal output
rlabel metal2 s 66534 109200 66590 110000 6 o[78]
port 363 nsew signal output
rlabel metal2 s 67362 109200 67418 110000 6 o[79]
port 364 nsew signal output
rlabel metal2 s 7746 109200 7802 110000 6 o[7]
port 365 nsew signal output
rlabel metal2 s 68190 109200 68246 110000 6 o[80]
port 366 nsew signal output
rlabel metal2 s 69018 109200 69074 110000 6 o[81]
port 367 nsew signal output
rlabel metal2 s 69846 109200 69902 110000 6 o[82]
port 368 nsew signal output
rlabel metal2 s 70674 109200 70730 110000 6 o[83]
port 369 nsew signal output
rlabel metal2 s 71502 109200 71558 110000 6 o[84]
port 370 nsew signal output
rlabel metal2 s 72330 109200 72386 110000 6 o[85]
port 371 nsew signal output
rlabel metal2 s 73158 109200 73214 110000 6 o[86]
port 372 nsew signal output
rlabel metal2 s 73986 109200 74042 110000 6 o[87]
port 373 nsew signal output
rlabel metal2 s 74814 109200 74870 110000 6 o[88]
port 374 nsew signal output
rlabel metal2 s 75642 109200 75698 110000 6 o[89]
port 375 nsew signal output
rlabel metal2 s 8574 109200 8630 110000 6 o[8]
port 376 nsew signal output
rlabel metal2 s 76470 109200 76526 110000 6 o[90]
port 377 nsew signal output
rlabel metal2 s 77298 109200 77354 110000 6 o[91]
port 378 nsew signal output
rlabel metal2 s 78126 109200 78182 110000 6 o[92]
port 379 nsew signal output
rlabel metal2 s 78954 109200 79010 110000 6 o[93]
port 380 nsew signal output
rlabel metal2 s 79782 109200 79838 110000 6 o[94]
port 381 nsew signal output
rlabel metal2 s 80610 109200 80666 110000 6 o[95]
port 382 nsew signal output
rlabel metal2 s 81438 109200 81494 110000 6 o[96]
port 383 nsew signal output
rlabel metal2 s 82266 109200 82322 110000 6 o[97]
port 384 nsew signal output
rlabel metal2 s 83094 109200 83150 110000 6 o[98]
port 385 nsew signal output
rlabel metal2 s 83922 109200 83978 110000 6 o[99]
port 386 nsew signal output
rlabel metal2 s 9402 109200 9458 110000 6 o[9]
port 387 nsew signal output
rlabel metal2 s 107934 109200 107990 110000 6 rst
port 388 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 110000 110000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 44622574
string GDS_FILE /scratch/mpw7/caravel_user_project/openlane/multiply_add_64x64/runs/22_12_05_18_26/results/signoff/multiply_add_64x64.magic.gds
string GDS_START 287814
<< end >>

